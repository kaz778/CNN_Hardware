////round(2^k)

////conv1.weight

//parameter filter_28_24 = 25'b00000_11101_11100_11110_11000;

////conv2.weight

//parameter filter_12_8_1 = 25'b11111_10000_10000_10001_10011;
//parameter filter_12_8_2 = 25'b10000_10000_10000_10111_11111;
//parameter filter_12_8_3 = 25'b10000_10000_11111_11110_00000;
//parameter filter_12_8_4 = 25'b00000_00000_00111_01110_01100;

////fc1.weight

//parameter fc_64_16_0 = 64'b11111_10000_01111_01001_11110_10110_00100_10101_01101_00100_00111_10000_0001;
//parameter fc_64_16_1 = 64'b01011_11101_10001_00000_11011_11111_10111_11100_11101_11000_00111_01011_1111;
//parameter fc_64_16_2 = 64'b10101_01010_01001_11101_11100_01100_00000_10110_01100_01111_00110_01101_0001;
//parameter fc_64_16_3 = 64'b01111_10011_01000_10111_00110_00000_11000_01001_10010_01101_11001_10110_0000;
//parameter fc_64_16_4 = 64'b00010_11111_01111_11101_00000_00010_11101_10001_01000_00000_11001_00110_0110;
//parameter fc_64_16_5 = 64'b11111_10010_00000_00001_00111_01101_00111_11101_10001_11010_00111_11101_1101;
//parameter fc_64_16_6 = 64'b11010_01100_10000_01001_00000_11001_00001_10011_00100_11011_10100_10000_0111;
//parameter fc_64_16_7 = 64'b11111_11001_10100_10111_00000_11011_00110_01001_11000_01000_11110_10011_0010;
//parameter fc_64_16_8 = 64'b01110_00100_10111_10110_10011_00011_00000_01111_10111_11100_01110_10000_1110;
//parameter fc_64_16_9 = 64'b10001_10001_00111_10111_01010_10011_01111_11101_11010_00010_01110_01011_0110;
//parameter fc_64_16_10 = 64'b00000_01011_10111_10011_00001_00011_11110_11110_11100_00111_01110_01100_1100;
//parameter fc_64_16_11 = 64'b01111_10110_00000_00011_10011_01110_10100_01011_00010_11100_00011_01100_1000;
//parameter fc_64_16_12 = 64'b00001_11011_10000_00000_10001_11011_10111_11100_10000_11110_00110_01111_1111;
//parameter fc_64_16_13 = 64'b00011_10110_01011_01101_01001_10110_01111_11101_10010_00000_00111_01110_1001;
//parameter fc_64_16_14 = 64'b10100_01101_00110_01010_11111_00000_00011_00111_11101_10011_11001_10111_1001;
//parameter fc_64_16_15 = 64'b11000_00010_11010_01000_00001_01111_11001_10011_10011_11111_10000_00000_1110;

////fc1.bias

//parameter fc_64_16_bias = 16'b10110_00000_11110_1;

////fc2.weight

//parameter fc_16_10_0 = 16'b01100_01100_00101_0;
//parameter fc_16_10_1 = 16'b11011_00010_01010_0;
//parameter fc_16_10_2 = 16'b11100_10000_01111_0;
//parameter fc_16_10_3 = 16'b11000_10111_11100_1;
//parameter fc_16_10_4 = 16'b10010_00011_10001_0;
//parameter fc_16_10_5 = 16'b01000_01010_11001_1;
//parameter fc_16_10_6 = 16'b10110_11110_01001_0;
//parameter fc_16_10_7 = 16'b01011_00101_10111_0;
//parameter fc_16_10_8 = 16'b00110_10000_11100_1;
//parameter fc_16_10_9 = 16'b10101_01001_10011_1;

////fc2.bias

//parameter fc_16_10_bias = 10'b00111_01010;



////round(2^k-1)

////conv1.weight

//parameter filter_28_24 = 25'b00000_10000_00001_00001_00111;

////conv2.weight

//parameter filter_12_8_1 = 25'b00000_00000_11111_11000_00000;
//parameter filter_12_8_2 = 25'b01110_00111_00001_00000_00000;
//parameter filter_12_8_3 = 25'b11000_10000_10010_00000_00000;
//parameter filter_12_8_4 = 25'b00000_10000_00000_11100_11110;

////fc1.weight

//parameter fc_64_16_0 = 64'b00001_10100_01010_00000_01101_01111_11001_11000_11011_10111_11010_10001_1000;
//parameter fc_64_16_1 = 64'b11001_11000_00111_01100_11001_10000_00000_11001_00110_01011_10001_00010_1111;
//parameter fc_64_16_2 = 64'b11101_10010_11111_01011_00110_00100_10110_11000_00011_00111_00011_11011_1110;
//parameter fc_64_16_3 = 64'b10110_01111_00000_01000_01000_01110_01111_01010_00100_11000_11111_10010_0000;
//parameter fc_64_16_4 = 64'b00010_11111_11101_11001_10000_10010_10000_01110_01001_10000_11010_11110_1001;
//parameter fc_64_16_5 = 64'b00010_00001_01110_00111_01110_11011_11011_10111_11101_10100_00000_00000_1000;
//parameter fc_64_16_6 = 64'b10111_11000_00000_01110_00101_11110_01110_10001_01110_01111_10101_00001_1000;
//parameter fc_64_16_7 = 64'b11100_00100_11111_10011_10010_10000_00110_01100_10001_00111_11001_10111_1110;
//parameter fc_64_16_8 = 64'b11101_01100_00000_00000_00001_00100_11100_00101_11110_00010_11101_10000_0000;
//parameter fc_64_16_9 = 64'b11100_00100_10000_00111_00011_00001_00011_01110_00100_01000_01001_10111_1110;
//parameter fc_64_16_10 = 64'b10010_00011_00011_11111_11110_01110_00111_11001_00110_01110_00010_01010_0111;
//parameter fc_64_16_11 = 64'b11000_00101_10001_11110_00110_01100_01110_01101_10011_10010_01111_10100_0010;
//parameter fc_64_16_12 = 64'b00000_00000_01011_10100_01001_11111_11001_10111_10010_01000_00000_00010_0110;
//parameter fc_64_16_13 = 64'b01000_01001_00011_10000_01111_11111_10101_01111_11010_00000_11001_00110_0111;
//parameter fc_64_16_14 = 64'b11010_01101_11000_00010_10111_11111_10101_11100_11010_10100_01010_10101_0100;
//parameter fc_64_16_15 = 64'b11110_00010_10101_10011_11111_11110_10000_10111_11010_00010_00000_01100_1111;

////fc1.bias

//parameter fc_64_16_bias = 16'b01010_11011_10100_0;

////fc2.weight

//parameter fc_16_10_0 = 16'b10111_10111_01101_0;
//parameter fc_16_10_1 = 16'b01010_11001_10100_0;
//parameter fc_16_10_2 = 16'b10011_01000_01000_0;
//parameter fc_16_10_3 = 16'b11101_00100_00000_0;
//parameter fc_16_10_4 = 16'b11100_11000_11111_1;
//parameter fc_16_10_5 = 16'b00101_10101_10000_1;
//parameter fc_16_10_6 = 16'b10011_11011_00011_1;
//parameter fc_16_10_7 = 16'b01110_01111_11001_0;
//parameter fc_16_10_8 = 16'b00011_10000_11011_0;
//parameter fc_16_10_9 = 16'b01000_00111_01111_1;

////fc2.bias

//parameter fc_16_10_bias = 10'b11000_01001;



//floor(2^k)

//conv1.weight

parameter filter_28_24 = 25'b01111_01111_11110_00000_00000;

//conv2.weight

parameter filter_12_8_1 = 25'b01000_01111_11111_00001_00000;
parameter filter_12_8_2 = 25'b11101_10000_10000_10001_00011;
parameter filter_12_8_3 = 25'b00111_01111_11100_00000_00000;
parameter filter_12_8_4 = 25'b01000_00000_01110_11110_11110;

//fc1.weight

parameter fc_64_16_0 = 64'b00010_01100_11111_11111_11100_11011_10011_10011_01001_01101_00110_01101_1100;
parameter fc_64_16_1 = 64'b00101_00000_01001_11111_11111_01100_00111_00110_00110_00100_11000_01100_1101;
parameter fc_64_16_2 = 64'b01101_11100_11000_01000_00011_00111_11000_01100_10110_11011_11100_10000_0010;
parameter fc_64_16_3 = 64'b01110_00111_11011_11110_11100_00000_00111_11111_00010_00111_01100_11101_1011;
parameter fc_64_16_4 = 64'b01110_00111_11110_01111_00000_00000_01011_10001_10011_10011_01111_10101_0001;
parameter fc_64_16_5 = 64'b01111_11100_00011_11000_00000_01100_10011_00110_10010_00011_11100_10100_1001;
parameter fc_64_16_6 = 64'b00011_11110_11100_00110_01111_11011_11001_11011_10010_01011_01011_00010_0000;
parameter fc_64_16_7 = 64'b00011_00100_11101_00111_01111_00010_11011_10011_00100_00101_10111_00111_0001;
parameter fc_64_16_8 = 64'b01000_11111_00010_00000_00000_11011_01000_01100_11111_11110_01100_11001_0000;
parameter fc_64_16_9 = 64'b11001_00000_01001_11010_01010_00100_10010_01001_00110_00011_01010_11111_1001;
parameter fc_64_16_10 = 64'b11011_11111_10111_10111_10110_00000_00111_11000_01001_00000_00001_01011_1111;
parameter fc_64_16_11 = 64'b00000_01000_01110_11110_01100_10011_01000_10110_00001_01111_00110_11001_0000;
parameter fc_64_16_12 = 64'b00110_00010_11100_01111_01100_00110_11001_10000_00101_10001_10101_10110_0010;
parameter fc_64_16_13 = 64'b00001_10000_01111_11111_11101_10010_10111_11100_00011_11100_00100_11111_0000;
parameter fc_64_16_14 = 64'b00110_01100_10000_01111_00101_11000_10011_10010_01100_00101_10100_01001_1111;
parameter fc_64_16_15 = 64'b11001_10100_01000_10001_10001_11000_00111_01010_01100_01110_11000_11001_1111;

//fc1.bias

parameter fc_64_16_bias = 16'b11000_00101_10101_1;

//fc2.weight

parameter fc_16_10_0 = 16'b11010_10010_01001_1;
parameter fc_16_10_1 = 16'b01000_01100_00100_1;
parameter fc_16_10_2 = 16'b01010_10001_10010_1;
parameter fc_16_10_3 = 16'b00011_00011_10000_1;
parameter fc_16_10_4 = 16'b10011_00111_01110_0;
parameter fc_16_10_5 = 16'b10011_11010_10001_0;
parameter fc_16_10_6 = 16'b11011_00100_11111_1;
parameter fc_16_10_7 = 16'b00100_11010_01010_1;
parameter fc_16_10_8 = 16'b01111_11101_00001_1;
parameter fc_16_10_9 = 16'b00101_10010_01110_0;

//fc2.bias

parameter fc_16_10_bias = 10'b10010_01010;
