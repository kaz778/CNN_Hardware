parameter data_0 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010010110_011111101_011001010_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111011_011111011_011111101_001101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011000101_011111011_011111011_011111101_001101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_010111110_011111011_011111011_011111011_011111101_010101001_001101101_000111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111011_011111011_011111011_011111011_011111101_011111011_011111011_011011100_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110110_011111111_011111101_011111101_011111101_011111101_011101010_011011110_011111101_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011011101_011111101_011111011_011111011_011111011_010010011_001001101_000111110_010000000_011111011_011111011_001101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011100111_011111011_011111101_011111011_011011100_010001001_000001010_000000000_000000000_000011111_011100110_011111011_011110011_001110001_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111011_011111011_011111101_010111100_000010100_000000000_000000000_000000000_000000000_000000000_001101101_011111011_011111101_011111011_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111011_011111011_011001001_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011001000_011111101_011111011_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011001010_011111111_011111101_010100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111011_011111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011111011_011111101_011111011_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011001_011111011_011111011_000000000_000000000_000000000_000000000_000000000_000000000_000010101_000111111_011100111_011111011_011111101_011100110_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011001_011111011_011111011_000000000_000000000_000000000_000000000_000000000_000000000_010010000_011111011_011111011_011111011_011011101_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011001_011111011_011111011_000000000_000000000_000000000_000000000_000000000_010110110_011011101_011111011_011111011_011111011_010110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011010_011111101_011111101_001001001_001001001_011100100_011111101_011111101_011111111_011111101_011111101_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011111011_011111011_011111101_011111011_011111011_011111011_011111011_011111101_011111011_011111011_011111011_010010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011100110_011111011_011111101_011111011_011111011_011111011_011111011_011111101_011100110_010111101_000100011_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111110_010001110_011111101_011111011_011111011_011111011_011111011_011111101_001101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_010101110_011111011_010101101_001000111_001001000_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_1 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_000000011_000101010_001110110_011000001_001110110_001110110_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_010110011_011110101_011101100_011110010_011111110_011111110_011111110_011111110_011110101_011101011_001010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010111_011111110_011111110_011111110_011010101_011000000_010110010_010110010_010110100_011111110_011111110_011110001_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011101011_011111110_011100010_001000000_000011100_000001100_000000000_000000000_000000010_010000000_011111100_011111111_010101101_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111000_011111110_011111101_001101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011111010_011111110_001001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011111110_010011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011101_011111110_010011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000010_011111110_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010110_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011011100_011101111_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111110_011111110_010101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010110_011101111_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010110_011000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_011011011_011000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111110_011000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111110_011010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111110_011000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011101110_011111110_001001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111110_011000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_010100101_011111110_011000011_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011110001_011000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_010100111_011111110_011100011_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010110_011010101_000010100_000000000_000000000_000000000_000000000_000000000_000101110_010011000_011001010_011111110_011111110_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010110_011111110_011001100_010110100_010110100_010110100_010110100_010110100_011101011_011111110_011111110_011101010_010011100_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_011001101_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111100_011101010_001111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011010010_011111110_011111110_011111110_011111110_011111110_010011001_001101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_2 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_001000010_010001010_011111111_011111101_010101001_010001010_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001111000_011100100_011111100_011111100_011111101_011111100_011111100_011111100_010011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101100_011111100_011111100_011111100_011111100_010111110_011111100_011111100_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011101001_011111100_011111100_011111100_001110100_000000101_010000111_011111100_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_010110010_011111101_011111100_011011101_000101011_000000010_000000000_000000101_000110110_011101000_011111100_011010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_011111101_011111111_011111001_001110011_000000000_000000000_000000000_000000000_000000000_010001000_011111011_011111111_010011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100110_011111100_011111101_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010001_011111101_011001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011011100_011111100_011111101_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_011111100_011111100_011000000_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011011111_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111010_011111100_011111100_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011111100_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111111_011111101_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111000_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011111100_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111000_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011110000_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111000_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010010_011111101_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_011101000_011111100_010011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100110_011101000_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_011111101_011110100_000110010_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011111101_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_010100100_011111101_001110001_000000000_000000000_000000000_000000000_000000000_001000010_011101100_011100111_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011011110_011110000_010000110_000000000_000000000_000100110_001011011_011101010_011111100_010001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_010110001_011110000_011001111_001100111_011101001_011111100_011111100_010110000_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_000110110_010110011_011111100_010001001_010001001_000110110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_3 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001010000_011000011_001010101_001010000_001010000_001010000_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011111101_011111101_011111101_011111101_011111101_011111101_010011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_000111110_000111000_000000000_000001001_011111101_011111101_011111101_011111101_011111101_011111101_011111011_011101101_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111101_011110001_001010011_000000100_010100001_011111101_011111101_011111101_011111101_011111101_011111101_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010001101_011111000_011111101_011111101_010010011_000000000_001001001_011010001_011111100_011111101_011111101_011111101_011111101_011111101_011010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010011_011111101_011111101_011111101_011111101_011000111_000100010_000000000_000000000_010100000_011111101_010001110_011000010_011111101_011111101_011110100_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010001000_011111010_011111101_011111101_011111101_011111101_011111101_001000101_000000000_000000000_000001111_000110100_000000101_000011011_011001001_011111101_011111101_010011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010000_011111101_011111101_011111101_011111101_011111101_011111101_011010001_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011111101_011111101_011000100_000100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111101_011111101_011111101_011111101_011111101_011101010_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101010_011111101_011111101_011111101_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011111101_011111101_011111101_011111101_010100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_011111101_011111101_011111101_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011111101_011111101_011111101_010101100_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_011111101_011111101_011111101_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011111101_011111101_011010010_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000101010_011100101_011110110_011111100_011111101_011111101_010011111_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011111101_011111101_011010001_000000000_000000000_000000000_000000000_000000000_001100011_010010101_011010010_011111101_011111101_011111101_011111101_011110010_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111101_011111101_011111101_011011010_000110101_000110101_000110101_010110100_011100100_011110100_011111101_011111101_011111101_011111101_011111101_011111101_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011000001_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010000_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011101010_011000001_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011010010_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011100101_001000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011100100_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111000_011101011_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100111_011010010_011111101_011111101_011111101_011111101_011111101_011111101_010111101_001110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_001101100_011111101_011111101_010110011_001001110_001001110_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_4 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011111111_011111110_011111111_011111110_011111110_011111110_010011101_010000010_001011000_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_001101100_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_010000001_011101110_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111000_011111101_011111000_010100111_011101011_011111101_011111101_011111101_011111101_001101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_010110010_011111101_010110110_000000000_000011011_010000110_011110111_011111101_011111101_011010111_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_010000010_011111101_011011110_000011011_000000000_000000000_000000000_010111010_011111101_011111101_011111101_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011111101_011111101_001111010_000000000_000000000_000000000_000000000_001000011_011110110_011111101_011111101_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110101_011111101_011000111_000011001_000000000_000000000_000000000_000000000_000000000_010111011_011111101_011111101_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_011100001_011110101_001000011_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111101_011111101_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010101_011111101_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111101_011111101_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011100100_011111101_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111101_011111101_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011111101_011111101_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111101_011111101_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011111101_011111101_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111101_011111101_001101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011111101_011111101_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111101_011011011_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011111101_011111101_011100110_000100000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111101_010011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011111101_011111101_011111101_011101001_001111000_000000000_001001010_001100100_001100100_011001000_011111000_011011001_000100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_010011111_011111101_011111101_011111101_011111001_011100110_011110111_011111101_011111101_011111101_011111101_001101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_001110110_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_000101001_011111101_011111101_011111101_011111101_011111101_011111101_011111101_001110111_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_000110011_001011000_011010110_010100101_001100011_000000101_000000101_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_5 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_000011101_000000100_001101000_011100101_011111101_010000001_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011111100_010110011_011111100_011111100_011111100_011111101_001111010_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011111100_011111101_011111100_010010100_000111000_011111101_011111100_010001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011110110_011111100_011111101_001100110_000000110_000000000_010011001_011111100_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101010_011111101_011111101_011111111_001010100_000000000_000000000_000001101_011001111_011111101_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_011111100_011110111_001000001_000000000_000000000_000000000_010101001_011111100_011010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_011111100_001100100_000000000_000000000_000000000_000000000_001010010_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011110011_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000111001_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011111101_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000111001_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111100_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000111001_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100101_011111100_011100000_010101000_000000000_000000000_000000000_000000000_000000000_000111001_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_010101000_000000000_000000000_000000000_000000000_000000000_000000000_001111000_011111101_010111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_001011101_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_000111000_000000000_000000000_000000000_000000000_000000000_000001010_011000101_011111100_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_010011100_000000000_000000000_000000000_000000000_000000000_010110011_011111100_010110001_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110011_011111101_010110010_000010000_000000000_000010011_001000010_010111111_011111110_011010001_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011101010_011111100_011010111_010101001_011100001_011111100_011111100_011010001_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000011_011111100_011111100_011111101_011111100_011111100_011010110_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_001000001_011110000_011111101_010110001_001100111_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_6 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101111_011011001_011101000_010000100_000111001_001011100_001011100_001011100_001011100_000101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_010011111_011111100_011111110_011111110_011111110_011111100_011111110_011111110_011111110_011111110_011111011_010001001_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011001101_011111110_011111110_011111110_011111110_011111110_011101010_011001000_010000101_010000101_011000101_011110010_011111110_010110010_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011100000_011111110_011100000_011001000_001111100_010001010_011001000_000100000_000000000_000000000_000000000_000000000_000100110_010110100_011111110_010000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011011111_011111110_011101111_000100001_000000100_000000000_000000000_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011101011_011110000_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001110111_011111110_011111001_001000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111110_011111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011111110_011111110_001100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_011111110_011111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010000_011111110_011101100_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_011111110_011111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111100_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001001_011111110_011111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011110100_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111110_011000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111110_001000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011110111_011111110_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111110_001001010_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001001100_011011110_011111110_011101000_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011111110_011111110_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_001110001_011000000_011111110_011111110_011001111_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_011011110_011111110_011111000_010111001_010000110_001100011_000111110_010000110_010000110_010000110_011001000_011110011_011111110_011111110_011101001_010001011_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_010100010_011111100_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111000_001111110_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_010101100_010111010_010111010_011010100_010111010_010111010_010111010_001111010_001011011_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_7 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111110_011111110_011111110_011111110_010000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011010_011111010_011111101_011111101_011111101_011111101_011111100_011111000_010100000_001110110_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011000_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011101000_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010000_011111011_011111101_011111101_011100000_000110000_000110001_010101010_011111101_011111101_011111101_011111101_011101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011111011_011111101_011111101_010110110_000010010_000000000_000000000_000000110_000110001_010101010_011111101_011111101_011111011_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011100001_011111101_011111101_011111101_000111101_000000000_000000000_000000000_000000000_000000000_000011010_011011101_011111101_011111101_011110101_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_011110101_011111101_011111101_011111101_010001001_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000101010_011011101_011111101_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111101_011111101_011111101_011100001_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011100_011111101_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111101_011111101_011111101_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011100_011111101_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010111_011111101_011111101_010110001_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011100_011111101_011111101_011011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111000_011111101_011111101_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011100_011111101_011111101_011110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011111101_011111101_001111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011100_011111101_011111101_011011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010000_011111101_011111101_010011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_010101110_011111101_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100000_011111101_011111101_010011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_010000110_011111101_011111101_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111101_011111101_010011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_001000011_011111101_011111101_011111101_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_011110110_011111101_011011000_000100001_000000000_000000000_000000000_000000000_000000111_000011011_010000110_011111101_011111101_011111101_011111011_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011110001_011111101_011111101_011011000_000101000_010000000_010010110_010010110_010101110_011111101_011111101_011111101_011111101_011111011_011010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101001_011110011_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100101_011111101_011111101_011111101_011111010_011111101_011111101_011011101_011010010_010011100_010110111_001110101_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100001_010001011_011101010_001010011_001111011_001111011_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_8 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011000011_011100100_001000000_001010010_010011100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011100000_011111101_011111110_011111001_011010100_011111101_011010000_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001001_011001011_011111101_011100011_011010000_011111101_001110000_011010101_011111101_011001101_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011111001_011111101_010100111_000101001_010010111_010110110_000010101_001100111_011110110_011111110_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111110_011111101_011001111_000100011_000000000_000000000_000000000_000000000_000000110_001001111_010111101_011101101_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_011111110_011111111_011111110_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101010_011111110_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011100000_011111101_011111110_010000010_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_010011000_011100000_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111101_011111101_010011111_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_011110111_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001100_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_011101000_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011111_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011110000_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111010_011111110_011100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011110011_000100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111010_011111101_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101010_011101001_011011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011111101_011111101_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110111_011111101_010101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011100111_011111101_001010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_011101010_011111101_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111110_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_010110101_011111110_010110101_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011010100_011111110_010101010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_010100111_011111110_011101010_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011111101_011111110_001100101_000001000_000000000_000000000_000000000_000110011_010011110_011111001_011101001_001101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_010001011_011111110_011111101_011011110_010110010_010000000_011011010_011101110_011111101_011100111_000110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_010010000_011100100_011111010_011111101_011111101_011111110_011111001_010111101_001010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111110_001001000_010101001_001101001_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_9 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101010_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_001100010_010011101_011111100_011101111_011010001_001010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_011011000_011111110_011111110_011111110_011111110_011111110_011111010_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_010111111_011111011_011000111_010001011_000111101_000111101_010101101_011111111_010001101_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_010111111_011111110_011110001_000000000_000000000_000000000_000000000_000010000_010101111_011111110_011010111_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011001111_011111110_011100010_001100001_000000000_000000000_000000000_000000000_000000000_000001100_010111101_011111110_011010101_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111100_010101000_011111110_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001010_011111110_011111110_011010110_001100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101011_011111110_011100110_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000001_001001010_011111001_011111110_011111101_010000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101010_011111100_011100100_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000001_011111110_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111110_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_010111110_011111110_011110111_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000001_011111110_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111110_011111110_011000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111110_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_011111001_011111110_011101100_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111110_001111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000101_011111110_011111110_001111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111110_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011111110_011111110_010111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_011101100_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011111110_011110110_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101011_011001011_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011001000_011111110_011110000_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100111_011010011_001101101_000111111_000111111_000111111_000111111_000011101_000111111_000011101_000111111_000111111_000111111_011000010_011011010_011111110_011111110_011101110_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_001101001_011110001_011111110_011111110_011111110_011010110_011111110_011010110_011111110_011111110_011111110_011111110_011111110_011110100_001110100_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000001_010110010_011101010_011101010_010111001_011010000_011101010_011101010_011101010_010100110_001100000_001100000_001001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_10 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011111110_001101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010111_011111100_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_011110100_010010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111110_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001010_011011111_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011111110_011011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011111110_011000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111110_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011101101_011001101_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111100_011111111_010100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101011_011111110_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011101000_011010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111000_011111110_010011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010111_011111110_010001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100100_011111110_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_011111011_011111110_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111110_011001101_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011010111_011111110_001111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_011000110_010110000_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_11 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001101_011111110_001101011_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011100011_011111110_011111110_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_011111110_011111110_010100101_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011001011_011111110_011111110_001001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_011111110_011111110_011111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011111110_011111110_010110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000100_011111110_011111000_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111010_011111110_011111110_011101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101111_011111110_011111110_010000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011111110_011101110_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111100_011111100_011111110_011011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011111110_011111110_010011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011111110_011101110_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011111100_011111110_011010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111110_011111110_010000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101001_011111110_011101010_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101111_011111110_011001100_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_011010011_011111110_011000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_010011110_011111110_010100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_010011101_001101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_12 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_13 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011010_011111101_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011001_011111100_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001000_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011001100_011111010_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011111001_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011111100_011110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001111_011111100_011110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111110_011111100_011110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100000_011111100_011110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100101_011111100_011111101_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_010111000_011111111_010101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111101_011100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111101_011100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111101_011100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111101_011100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010101_011111101_011101011_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001001_011111101_011111100_001100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111101_011111100_001100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111101_011111100_001100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011000011_011110001_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_14 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011000001_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011111101_010000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111110_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111101_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011111110_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011000_011111101_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011000_011111100_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011111101_011010110_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011010100_011111101_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011111110_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111101_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111110_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111101_011000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111110_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111101_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011111111_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101101_011111101_000111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_15 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011011010_011010001_000111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_010111101_011111100_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_011010111_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_011111101_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_011111101_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011111101_011111110_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111100_011111101_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111011_011111001_011111101_011010010_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010100_011111111_011111101_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100111_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010100_011111111_011111101_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000011_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101010_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101010_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_011010001_010110110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_16 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011011110_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011011111_011111110_001111111_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011111110_011111110_011111110_010101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110101_011111110_011111110_011111110_010101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110101_011111110_011111110_011111110_010011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110101_011111110_011111110_011110011_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011100110_011111110_011111110_010110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011111110_011111110_011111110_010011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011000000_011111110_011111110_011111110_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011111110_011111110_011111110_011111110_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011111110_011111110_011111110_011101100_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011111110_011111110_011111110_010111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011111110_011111110_011111110_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011111110_011111110_011001010_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011010111_011111110_011110110_001100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011011111_011111110_011111110_010111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011010000_011111110_011111110_010111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011010111_011111110_011111110_010111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011011001_011111110_011111110_010111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011111111_011111111_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_17 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100001_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011001_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000101_011100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011101010_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_001010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011111111_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011111110_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011101001_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_011100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100111_011010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100111_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011101001_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011111101_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_18 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010111_011111101_010100111_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_011011110_011111100_011111100_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_011111100_011111100_010111011_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111100_011111100_011111100_001011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_011111000_011111100_011111100_010001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000001_011111100_011111100_011100101_000100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_011111100_011111100_011111100_011010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011101011_011111100_011111100_011100010_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111100_011111100_011111101_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_011000011_011111100_011111101_011001001_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111100_011111101_011111111_011111101_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011110_011111100_011111101_011111100_001111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011111100_011111101_011111100_011000000_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_011010100_011111101_011111100_011111100_001110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101111_011111101_011111100_011111100_011000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011111101_011111100_011111100_011101110_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001000_011111100_011111100_011111100_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111101_011111100_011111100_011111100_011000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011111100_011111100_011111100_001110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001101110_011101001_011110011_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_19 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001101_011111110_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011111101_011011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_001100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011110111_001001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011111110_011100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111110_010000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011110010_011111110_001101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100100_011111100_011110011_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011111101_001111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011101000_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111101_011101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110010_011111101_001101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011010_011111101_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011010_010101010_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011100110_010010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011111101_010010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011011101_010010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100000_011000100_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_20 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_001111101_010101011_011111111_011111111_010010110_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111101_011111101_011111101_011111101_011111101_011111101_011011010_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111101_011111101_011111101_011010101_010001110_010110000_011111101_011111101_001111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110100_011111010_011111101_011010010_000100000_000001100_000000000_000000110_011001110_011111101_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001101_011111011_011010010_000011001_000000000_000000000_000000000_001111010_011111000_011111101_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_000010010_000000000_000000000_000000000_000000000_011010001_011111101_011111101_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110101_011110111_011111101_011000110_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001100_011110111_011111101_011100111_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111101_011111101_010010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110000_011110110_011111101_010011111_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_011101010_011111101_011101001_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_011111101_011111101_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011111000_011111101_010111101_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011001000_011111101_011111101_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011111101_011111101_010101101_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111000_011111101_011111101_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111000_011111101_011111101_000101011_000010100_000010100_000010100_000010100_000000101_000000000_000000101_000010100_000010100_000100101_010010110_010010110_010010110_010010011_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111000_011111101_011111101_011111101_011111101_011111101_011111101_011111101_010101000_010001111_010100110_011111101_011111101_011111101_011111101_011111101_011111101_011111101_001111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101110_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111001_011110111_011110111_010101001_001110101_001110101_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_001111011_001111011_001111011_010100110_011111101_011111101_011111101_010011011_001111011_001111011_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_21 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_001111101_010111111_011011010_011111111_011111110_011111110_011110001_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001100_011111001_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111010_011101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011110001_011111011_011111101_011100001_010001110_000110001_000001100_000001100_000001100_001101001_011111101_011111101_001101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011100001_011111101_010100111_001110001_000001110_000000000_000000000_000000000_000000000_000000000_000010000_011010011_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_011101110_011111101_010101010_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010110_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111011_011011010_000110000_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010110_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110000_011111101_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010111000_011110010_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_000101101_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_011111101_011110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011101010_011111000_001101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_010011101_011111101_010000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010111101_011111101_011001011_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010011100_011111101_011110110_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010011100_011111101_011001010_001000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010011100_011111101_011100010_001000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_000100001_000100001_010001100_010100011_010111010_011111101_011100010_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_001010001_011110100_011111101_011111101_011111101_011111101_011111101_011111101_011111101_010111010_001000110_000010111_000000000_000000000_000010110_010011100_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010000_011000011_011111101_011111101_011111101_011111101_011111101_011111000_011101010_010100110_011111000_011111101_011111101_011110000_010010110_001001001_010010000_001101000_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011111000_011111101_011111101_011111101_011111101_011111101_011110010_001101001_000000000_000000000_001101011_011110010_011111101_011111101_011111101_011110101_010100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011111010_011111101_011111101_011111101_011110111_010000111_000010101_000000000_000000000_000000000_000000000_000010101_001110101_010110111_010110111_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_001111011_010110000_010000111_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_22 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_010101010_011111110_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_010111111_011110101_011111110_011111110_010101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001000110_011110010_011111110_011101011_011101001_011111110_010110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_010111000_011111110_011110011_001100011_000011011_001101110_011111110_010110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011001101_011110111_001100010_000011010_000000000_000000000_001101110_011111110_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_001101000_000010100_000000000_000000000_000000000_000000000_001101110_011111110_000100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011010110_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011001000_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011100111_010010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011110100_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_011001001_010000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100100_011100010_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_001111010_011001101_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_001010100_011011000_011111010_010010000_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011001111_011100100_000100101_000000000_000000000_000000000_000000000_000010100_010001000_011101110_011111110_011100100_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011111110_001000010_000000000_000000000_000000000_000110101_010111110_011111110_011111110_011000101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011100111_010110110_000000000_000100000_001100101_010111000_011111001_011101111_010110011_001100000_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111110_001100011_010000000_011101000_011111110_011111011_010111001_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_011011101_011111110_011111110_011111110_011111110_011000000_001000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011111110_011111110_010111100_001101001_001001000_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_23 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_001100110_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011010110_011111101_010100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011101000_011011111_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011110100_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011110011_010100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011111101_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011101001_011010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010101101_011100000_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111100_010100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011111110_011000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011001011_011101001_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111101_001100110_000000000_000011111_000110011_000110011_000110011_001110001_001110000_001110001_010011000_010000100_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011111101_011111100_011011111_011001011_011101001_011111100_011111101_011111100_011111101_011111100_011111101_011111100_011111101_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_000110011_010101101_011111101_011111110_011111101_011111110_011010101_001100110_001100110_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011010101_011111100_011111101_011111100_011000000_001101111_000110010_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101101_011111101_011111111_011111101_011100000_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_011111101_010000010_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_001100110_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_24 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001100_010101110_011100010_011111111_010111001_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011110_001010011_001000100_001001010_010111010_011110011_001111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_000001011_000000000_000000000_000000111_001110010_011110010_001100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_001110010_011011110_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011011011_010100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_011011111_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011111001_001010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110110_010100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011010_010100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_011110001_010100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000001_011111110_001100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000001_011111110_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_001001111_001100110_000010100_000000000_000000000_010100101_010110101_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_010011111_011110010_011110110_011110110_011110010_001110111_000111011_011111101_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111011_011011111_000100011_000000000_000000101_001110100_011110011_011111110_011001111_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011110011_001100111_000000000_000000000_000000000_000000000_001010001_011111110_011011010_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011111110_000100000_000000000_000000000_000000000_001001110_011110100_011010110_011100010_011001000_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111110_000110010_000000000_000111000_001011101_011110101_011010110_000011110_000101010_011100011_011001010_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_011000000_011110001_011100110_011111101_011111110_010100111_000011101_000000000_000000000_000101000_010000110_011110100_010111000_001000101_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_010001001_010101101_001011110_000001100_000000011_000000000_000000000_000000000_000000000_000000001_001100110_011010001_011110000_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_25 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101111_010001000_011110001_011111110_011111110_011111110_011111110_011111110_011111111_011001010_010000010_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100001_011100100_011111101_011111101_011111101_011111101_011100111_010000111_010111111_011011010_011101010_011111101_011000011_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011110000_011111101_011111101_011111100_010111101_000011111_000000000_000000000_000000000_000100101_010010001_011111101_010110010_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_010110110_010110110_001000100_000000000_000000000_000000000_000000000_000000000_000000000_000000011_010001101_011111101_010011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_010110110_011110001_001010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110101_011111101_010101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_011111101_010101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_011111101_010101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011111101_010101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100110_011111101_001011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011000000_011001011_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001110010_011111101_010111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_011111101_011111101_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000110110_010000010_000010001_000000110_000000000_000000000_000000000_000000000_000000110_010111101_011111101_010010010_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_010110001_011111101_011111101_011111101_011000010_010010100_001111001_000000111_000000000_001111111_011111101_011101100_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_010111000_011111101_011010111_001100110_011001001_011010010_011111101_011111101_010111010_010100110_011110110_011111011_001111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011111101_011001010_000001101_000000000_000000000_000000111_001011010_011101010_011111101_011111101_011111101_011110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011111101_011101111_001101001_000001010_000000000_000101111_010011101_011101110_011111101_011111101_011111101_011111011_010000100_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_010101110_011111101_011111101_011011111_011011011_011101110_011111101_011111101_011011111_000110110_001011000_011111011_011111101_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000110010_011101000_011111101_011111101_011111101_011101010_001101100_000001100_000000000_000000000_001010011_011111101_011111010_001111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_26 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000100101_010000000_010001100_010001100_010001100_000111010_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101111_001110110_011000010_011111101_011111101_011111101_011111101_011111101_011111101_011010111_001010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011000110_011111101_011100101_010011011_000100001_000010100_000010100_000101010_001111100_011111011_011110111_010100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011101100_011110011_001101001_000000110_000000000_000000000_000000000_000000000_000000000_000000000_001101001_011111101_011110100_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011110010_011111101_001111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_011000111_011111101_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111101_001110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000000_011111101_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100111_001000000_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011110100_011100011_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111111_011111101_010001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111000_011111101_010001110_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_011111101_011010101_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111000_011100110_010110111_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_010100000_011111010_010110100_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000010_011111101_011001111_001001111_000010000_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_010011010_011111010_011111101_011111101_011111101_011101001_011101011_011011111_011100100_011100100_011100100_011001001_010000001_011101010_011110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_011111101_010000010_001010011_001010011_001010011_001010011_001000101_010001101_010001111_010011010_001011011_011010110_010001111_011100101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000100100_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_000000000_000010111_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_27 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_000010010_000010010_000110111_010001001_011000000_010000011_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_001011111_010100100_011111110_011111110_011111110_011111110_011111110_011111110_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_010010111_011001111_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111110_011111110_011111110_011111110_011111110_011010001_010011011_001000001_001000001_010010100_011111110_011110111_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_011101110_011111110_010100110_000101111_000010010_000000000_000000000_000000000_001110010_011111110_011111110_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_000011101_000000010_000000000_000000000_000000000_000000000_000000000_001110010_011111110_011111110_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011111010_011111110_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011111110_011111110_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111100_011111110_011111010_001001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_011111000_011111110_011100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111011_011111110_011111011_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011100101_011111110_011110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011010011_011111110_011111110_011110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_000101110_011100100_011111010_011111010_011111010_011111010_011111011_011111110_011111110_011111110_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_011111110_011111110_011111110_011111110_011111110_011111110_011111111_011111110_011111110_011111110_010010001_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_011100010_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011110100_001010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011101111_001100010_010101010_011011010_011111110_011111110_011110001_010011010_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011111110_011111110_011111110_011111110_011111110_011111110_010110110_000101001_000000000_000000000_000011000_001110010_011011100_011111110_011111110_010101110_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011111110_011111110_011111110_011111110_011111100_001010111_000001101_000000000_000000000_000000000_000000000_000000000_000010101_000111001_010110011_011111110_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011011000_011111110_011111110_010010101_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_010000111_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_28 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_001011110_010001001_010001001_011000000_010001001_010000011_000010010_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_000100100_010010011_000111001_011111110_011111110_011111110_011000111_011101111_011010101_010111110_011101100_001111101_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_000110110_010110011_011111110_011111110_011111110_011001001_001101111_010010001_001100110_000101110_000000000_000111110_011100010_010111000_010010110_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011111110_011111110_011111110_011111101_010101100_000011000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011101101_011111110_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011111110_011111110_011011001_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111110_011010101_011111110_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_001110110_000110011_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_010100001_011000111_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011100110_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001010100_011111110_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011111110_011111110_001001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011100100_011111110_011111110_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011111110_011111110_011111110_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101111_001100000_001100000_001100000_001100000_000010000_000000000_000000000_010010100_011111110_011111110_010001100_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_011011010_011110011_011111110_011111110_011111110_011111110_011101011_011101000_001111001_011110101_011111110_011000011_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011011100_011111110_011111110_011110000_001111100_001111100_001000101_000100001_000000101_000111111_011111100_011111110_011111110_010111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011111110_011111110_011000000_000000101_000000000_000000000_000000000_000000000_000001100_010111001_011111110_011111111_011111110_010111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_010111001_011111110_011101110_001000001_000000000_000000000_000000000_000000000_001001001_011000111_011111110_011010000_011001111_011101110_011101000_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011100011_011111110_011111110_001010000_000000000_000000000_000000000_000000000_001001010_011101110_011111110_010101101_000000010_000000000_001111100_011101100_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_011111110_011111110_011111110_000101111_000000000_000101001_001010100_010011110_011101111_011111110_001010101_000011110_000000000_000000000_000000000_001000101_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001111010_011111110_011111110_010111000_010010111_011101101_011000100_010000000_001011011_000100011_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001001001_001101010_011101001_010010101_010111100_000001001_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_29 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_010100100_011111110_011000101_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010101_010001101_010110011_011110010_010110100_011011111_011111110_011000100_001111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011001000_011111110_011111111_011111111_011111110_011101101_011101100_011101110_011110101_011111001_010100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011100110_011111110_011111110_011111110_011001111_001010111_000011010_000011001_000011011_000110001_011101111_011010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011100001_011111110_011111110_011111000_010000000_000000111_000000000_000000000_000000000_000000000_001000100_011111110_010111010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_011000001_011111110_011111110_011111110_001010010_000000000_000000000_000000000_000000000_000000000_000000000_001000111_011111110_011101111_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011111110_011111110_011111000_001010000_000000010_000000000_000000000_000000000_000000000_000000000_000000000_010011101_011111110_011010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011111110_011111110_010100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011011000_011111110_001111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_001001010_010010101_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111110_011011111_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000001_010111001_011111110_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_000100000_001011010_001111100_011111110_011111110_001100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_010101110_011101010_011111110_011111110_011111110_011100010_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010101_011111010_011111110_011111110_011111110_011111110_011111110_010111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111101_011111110_011111110_011111110_011111110_011111110_011111110_011101000_000101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011111100_011111110_011011111_011111110_011111110_011111110_011001100_001011111_011111100_011000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011111110_011111110_011111110_011111110_011111110_011100001_000011111_000000000_011110110_011100111_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011111110_011111110_011111110_011111110_010100111_000010101_000000000_000000000_011110110_011111110_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_011010000_011111110_011111000_010000101_000001001_000000000_000000000_000000000_010101110_011111110_010011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_010010110_000110110_000000000_000000000_000000000_000000000_000000000_010010100_011111001_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_001000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_30 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_000101001_010010010_010010010_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_010000001_011111101_011111101_011111101_011111010_010100011_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000101_011111101_011111101_011111101_011111101_011111101_011111101_011100101_001000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100101_011111101_011111100_010010001_001100110_001101011_011101101_011111101_011110111_010000000_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110101_011111101_010100111_000000000_000000000_000000000_000111101_011101011_011111101_011111101_010100011_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111101_000101011_000000000_000000000_000000000_000000000_000111010_011000001_011111101_011111101_010100100_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111011_011111101_000100000_000000000_000000000_000000000_000000000_000000000_000110111_011101100_011111101_011111101_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011111101_000100000_000000000_001100100_010111110_001010111_001010111_001010111_010010011_011111101_011111101_001111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011110_011111101_001001110_000101000_011111000_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011011111_001010100_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_001011100_000001100_000100011_011110000_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011110100_001011001_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_010100001_010110011_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011010001_000101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_000010000_000010000_000100111_000100110_000010000_000010000_010010001_011110011_011111101_011111101_010111001_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111010_011010001_011111101_011111101_010110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001101_011011101_011110111_001001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011011011_011111101_011110000_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011010_011110111_011111101_011111100_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_011111011_011111101_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011111101_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111100_011111101_010010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_010111100_011111101_011011101_010011110_000100110_000000000_000000000_000000000_000000000_001101111_011010011_011110110_011111101_011111101_010010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_011011101_011110110_011111101_011111011_011111001_011111001_011111001_011111001_011111101_011111101_011111101_011111101_011001000_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_010110111_011100100_011111101_011111101_011111101_011111101_011111101_011111101_011000011_001111100_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_000100101_010001010_001001010_001111110_001011000_000100101_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_31 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_001110001_011000001_011111110_011111101_011111110_011111101_011111110_010101100_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110111_011111101_011111100_011111101_011111100_011111101_011111100_011111101_011111100_011110011_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011111111_011101001_010110111_001100110_011001011_011001011_011101010_011111101_011111110_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_010010111_000110010_000000000_000000000_000000000_000101001_011000001_011111100_011111101_001101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_011010101_011111110_011111101_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011010101_011111100_011111101_011111100_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111101_011111110_011111101_011111110_010010111_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011010100_011111101_011111100_011111101_011101000_011011111_001111010_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011011111_011111110_011111101_011111110_011111101_011111110_001000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_000110010_010000011_011010101_011111100_011111101_011000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_010100010_011111110_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011001011_011111101_011111100_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111101_011111110_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_010001110_011111101_011111100_011101001_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011010110_011111101_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011110011_011111101_011111100_010101100_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010101101_010101101_011111101_011111111_011111101_011100000_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111100_011111101_011111100_011111101_010101011_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011001_011111101_011110100_011001011_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011000000_001111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_32 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111110_011111110_011111110_011111110_011011001_001110110_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110010_011110111_011111101_011111101_011111101_011111101_011111101_011111101_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011110100_011111101_011010000_010110001_010110001_000110111_001100011_011111101_011111001_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_010100101_010110011_000011001_000000000_000000000_000000000_001000101_011111101_011111101_001101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_011111101_011111001_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_010011001_011111101_010001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011110000_011111101_011111101_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_001101111_011110111_011111101_011111101_011100011_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011100100_011111101_011111101_011111101_011111101_011111101_011011101_001011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111100_011001110_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011001101_011001101_011001101_001010010_001000100_001000100_010111100_011111101_011111101_011100010_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111010_010100111_011111101_011111101_011100000_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_010110000_011111101_011111101_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101101_011111101_011011101_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101000_011111101_011111101_001001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011100011_011111101_011111101_001001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_000111111_010001100_011100010_011111101_011111101_011101110_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_000101010_010011001_011000001_011111101_011111101_011111101_011111101_011011001_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_000011101_010011110_011111011_011111101_011111101_011111101_011111101_011111101_011101000_001100110_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_001110100_010111010_011111101_011111101_011111101_011100011_001110100_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_33 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_010010111_011111111_011111110_010100011_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011010011_011111101_011111101_011111101_011111101_001000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011110001_010011000_010000111_011111000_011111101_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_001010100_000000000_000000000_010100010_011110111_011000000_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011000010_011111101_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111000_011111101_011111101_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011111101_011010000_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110100_011111101_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011101000_011111101_011001000_000111000_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011111101_011111101_011111101_011111101_010011111_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_010111001_011101011_011111101_011111101_011111101_010111110_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_001011001_011001001_011111101_011111101_011001110_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011010110_011111101_011111101_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001101_011111101_011111101_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_010000001_011110110_011111101_011011011_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001010_011001010_011111101_011111101_011011011_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100001_011100110_011110111_011111101_011111101_010101000_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100000_011111000_011111101_011111101_011111101_010000001_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100111_011111101_011111101_011111101_010000010_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101011_011111101_011100010_000100110_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_34 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_000111100_000111100_010000011_011010001_011010001_011010001_011010001_011010001_011010001_011010011_010101110_000111100_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001010_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011010011_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011111101_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_010110010_010110010_010110010_010110010_010110010_001100011_000011101_000011101_000011101_001011011_011110000_011111101_011111101_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_011110000_011111101_011111101_010100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_010000110_011111110_011111101_011111101_011111101_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_001011010_001011010_011101000_011110010_011111101_011111110_011111101_011111101_011111101_001101101_001010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_011010100_011111101_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011111101_011111101_011110110_001110100_000101110_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111000_011111101_011111101_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011111101_011111101_011111101_011111101_011111101_010010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111110_011111110_011111110_010011011_001111100_000000000_000000000_000000000_000000000_001001000_010010101_011100000_011111110_011111111_011111110_001101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_000101100_000101100_000101100_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_011100001_011111101_011111101_010001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_011110100_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011110110_011111101_010110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_011110001_010010001_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011110000_011111101_011111101_001101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_011111101_011111101_010110111_010110011_010110011_001110111_001000010_010110011_010110011_010110011_011101000_011111101_011110010_011000100_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011010110_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011111101_011111101_011111101_011111101_010100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_001011110_010100011_010110011_011001000_011111111_011111101_011111101_011111101_011100010_010100011_010100011_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_000011000_000111011_001011111_001101111_000111011_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_35 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011000000_001010111_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_011111101_010101010_000101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101111_011111001_011111101_011111100_011101001_001100101_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110011_011100011_011111100_011111100_011111100_010001010_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010111_001110000_010010011_011111100_011111100_010010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010000100_011110111_011111111_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110000_011111101_011000100_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111101_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010000100_011110110_011111101_010110110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011111101_011100011_010010100_010000011_001111011_011001001_011111101_011111101_011010100_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011111100_011111100_011111100_011111101_011111100_011111100_011100111_001111100_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_001001010_001111110_011010110_011101100_011111100_011111100_010010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_010001100_011111100_011100111_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011110100_011111100_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111100_000111110_000000000_000000000_000000000_000000000_000000000_000110010_011110101_011111101_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011110010_000011011_000000000_000000000_000000000_000100100_010010010_011010011_011111100_011111100_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_010110000_011111100_000010110_000010110_000011111_001111111_011011111_011111101_011111100_011110010_010000110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011111100_011111100_011111101_011111100_011111100_011111100_011111100_010111110_001101110_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_010110110_011111100_011111101_011111100_010011011_010010011_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_36 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_010000000_010000000_010000000_011111111_010000000_011111111_010111111_010000000_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_011111111_010111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_010000000_010000000_010000000_010000000_001000000_000000000_010000000_010111111_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_010000000_010000000_010111111_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_011111111_011111111_011111111_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_011111111_011111111_011111111_011111111_011111111_010111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_011111111_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_010111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_010000000_010000000_010000000_010000000_011111111_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_011111111_011111111_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_010111111_000000000_001000000_011111111_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_010111111_011111111_011111111_010111111_011111111_011111111_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_011111111_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_011111111_011111111_011111111_010000000_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_37 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_010101111_011100110_011111110_010000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011101100_011010001_011110101_011111110_011110010_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011101100_011001110_000110101_000100001_010010011_011111110_010010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110101_011011010_000001000_000000000_000000000_000100000_011110010_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_001101001_000000010_000000000_000000000_000100000_011101100_001001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_010100000_011011110_001010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011010111_011111110_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111110_011011001_011111110_010101101_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_010001111_011111010_011111110_011110101_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000011_011111110_011111110_011111110_011111110_011000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_011100000_011101111_010100100_011100101_010010111_010101111_001111110_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011100100_011111110_010101010_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010010100_011111110_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011011100_010110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111000_011101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111110_010011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_000001010_000000000_000000000_000000000_000000000_000000000_000000100_001010111_011001111_011111110_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_010100010_001111000_000000000_000000000_000000000_000000000_000000011_010010100_011111110_011111110_010101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011110101_011010000_000100100_000001100_000011000_001011001_011100001_011111110_011111110_011000110_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111101_011111111_011110111_011110001_011110100_011111110_011111111_011101010_001010000_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_38 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_010011100_011111101_011111101_011111111_011111101_011111101_011111101_010100101_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110000_011101101_011111100_011111100_011111100_011111101_011111100_011111100_011111100_011111100_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011100111_011100111_010100000_000100110_000010101_000010101_000101000_011111100_011111100_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_011111100_011111100_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011011111_011111100_011010000_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_010011101_011111101_011110011_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_010110111_011111100_011111100_011101101_001100110_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_001111111_011011111_011111101_011111100_011111100_011111100_011111100_011110010_010011001_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011001_011111100_011111100_011011000_010011001_001010100_010011010_011010111_011111101_011111100_011001010_000010101_000000000_000000000_000000000_000000000_000101011_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100100_011111100_010100100_000010010_000000000_000000000_000000000_000010010_001111010_011111100_011111100_011100001_000100011_000000000_000000000_001101011_010001101_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011100000_011111101_001111010_001101001_011100011_011011111_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011111100_011111100_011111101_010111101_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_001010101_011111100_011111100_010100001_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011000101_011111100_011111100_011111100_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011001_011101100_011111100_011111100_011111100_011111100_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_001000101_011101100_011010100_001001100_011110101_011111101_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100101_011111100_011011001_000101001_010111001_011111100_011111100_001000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011101010_011111100_001110000_011000000_011111100_011111011_010000110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011111100_011111100_011111100_011111101_011111100_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011111100_011111100_011111100_010111111_001110000_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_39 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_001110011_011000100_011111110_011111110_011111110_010011100_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000001_011001011_011111101_011111101_011111011_011111000_011111101_011111101_010011111_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_010001001_011111001_011111101_011110001_010010011_001000100_000101001_001110101_011110110_011111101_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011111101_011110010_010011101_000011101_000000000_000000000_000000010_001110011_011111010_011110111_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_010010001_000100100_000000000_000000000_000000000_000000000_000101101_011111101_011111101_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_001101111_010011001_011110000_011111101_011011011_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011111101_011111101_011111101_011100110_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010100_011101111_011111000_011111101_011111101_011111101_011111010_001100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101111_011111101_011111101_011111100_010110101_011111101_011111101_011111000_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000101100_000000100_000000100_000000001_000110010_010111000_011111101_011111100_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011100100_011111101_001111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111110_011111101_011011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000010_011111101_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101100_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100000_011111101_001111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011101100_010100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_001111000_011111010_011111101_001000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000001_011111101_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101111_011111101_011111101_010100101_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011101011_010110010_000000000_000000000_000000000_000000000_000000000_000010001_010011110_011110011_011111101_011001011_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011011_011101011_010001010_001011010_001011010_001011011_010010101_011011000_011111101_011111000_010100011_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111101_011111101_011111101_011111101_011111110_011111101_011101011_010010010_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_001111011_010100101_011111101_011000110_010011001_010000110_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_40 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010100_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_011000011_011100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100000_011010010_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_011111100_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_011101100_011011001_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000000_011111100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101000_011110111_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_011111111_011111101_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011110010_011010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111101_010111101_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011101000_011111010_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011100001_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011111100_011010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011111100_010100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_010100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011001100_011010001_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011111101_011111101_001101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111100_011000111_001010101_001010101_001010101_001010101_010000001_010100100_011000011_011111100_011111100_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_010101010_011110101_011111100_011111100_011111100_011111100_011101000_011100111_011111011_011111100_011111100_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_001010100_001010100_001010100_001010100_000000000_000000000_010100001_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111111_011111100_011111100_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111111_011111100_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011111100_011110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101000_011101100_001101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110011_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_41 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011000000_010000110_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_001001101_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011101011_011111010_010101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011011100_011110001_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_010111101_011111101_010010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001011_011111101_001100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_011111101_011111101_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011111110_010101101_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_010011001_011111101_001100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011100111_011111110_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011111111_011001100_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101000_011111110_010011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111101_010110010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010000011_011101101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111101_011111101_010111111_010101111_001000110_001000110_001000110_001000110_010000101_011000101_011111101_011111101_010101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011100100_011111101_011111101_011111110_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011011011_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_001000001_010001001_011111110_011101000_010001001_010001001_010001001_000101100_011111101_011111101_010100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011111110_011001110_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100000_011111101_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011111110_011110001_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011110_011111110_010100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100111_011110100_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101000_011111110_011101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010000_011111101_010011101_000000000_000001101_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010000_011111101_010011010_001011011_011001100_010100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010000_011111101_011111110_011111101_010011010_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_010111110_010000000_000010111_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_42 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101000_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_011101010_001111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111110_001111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_010110010_000011111_000000000_000000000_000000000_000000000_000000000_000110011_011111110_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011110_011111110_001010011_000000000_000000000_000000000_000000000_000000000_001010111_011111110_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100000_011111110_000111000_000000000_000000000_000000000_000000000_000000000_010111101_011101110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011100011_010101000_000000010_000000000_000000000_000000000_000000000_000000000_011000010_011101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011111110_001110010_000000000_000000000_000000000_000000000_000000000_000010000_011101011_010100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110011_011111110_000110010_000000000_000000000_000000000_000000000_000000000_001100111_011111110_001101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011011101_011101100_001001011_010011100_010110100_010111110_011111100_011111100_011111101_011111110_001110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011111110_011111110_011111110_011111100_011010011_010110011_010110011_010110011_011110110_011111110_011110111_001011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011011001_011101111_001110101_000010110_000000000_000000000_000000000_000000000_011100010_011111110_011110010_011000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_000010010_000000000_000000000_000000000_000000000_000000000_000011011_011110011_011001111_000101110_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111110_010000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111110_001000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111110_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111110_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101110_011111111_001100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111011_011111110_001010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110011_010110000_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_43 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011110011_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_010111010_011101100_000010101_000000000_000000000_000000000_010000110_001010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011010101_000011010_000000000_000000000_000000000_000000000_010000001_010101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_001111000_000000000_000000000_000000000_000000000_000000000_001011011_011010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011101010_001110000_000000000_000000000_000000000_000000000_000000000_001011011_011110010_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011011110_000010101_000000000_000000000_000000000_000000000_000000000_010101010_011110100_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_011110000_001111100_000000000_000000000_000000000_000000000_000000000_000101000_011111001_010001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001111111_011110001_000010010_000000000_000000000_000000000_000000000_000000000_000001111_011100110_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_011111110_010110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010111111_011101001_010001000_001100101_000010100_000000000_000000000_000000000_000000000_001110001_011010111_000011111_000011111_000011111_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_001011001_010000000_011000010_011011010_011010010_011010010_011010011_011010010_011100010_011111110_011111110_011001100_001111000_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_000001111_000100101_001011010_001011010_011000100_011110001_000100010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_011101001_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_010001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_010111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_011101001_000100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011111110_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_011010001_011011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101011_010100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_44 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011101_001110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111110_010010100_000000000_000000000_000000000_000000000_000010110_011100110_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101000_011111110_001110011_000000000_000000000_000000000_000000000_000011000_011111101_010111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011101010_011111110_001010001_000000000_000000000_000000000_000000000_001011011_011111101_010111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011011101_011111110_010100000_000000000_000000000_000000000_000000000_000000000_010001101_011111110_001111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011111101_011111101_001001100_000000000_000000000_000000000_000000000_000000000_011001111_011111101_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011101000_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_011001111_011111101_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100101_011111101_011001010_000010011_000000000_000000000_000000000_000000000_000000000_000100010_011110000_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_010101010_011111110_011111110_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000101111_011111110_011111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011111101_011111110_011111101_011101010_010100011_000101111_000101111_000011010_000000000_000000000_010000010_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011110110_011111110_011111101_011111101_011111101_011111110_011111101_011101000_010101110_011010000_011101000_011111101_010110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_010100001_011010011_011011011_011011011_011111110_011111101_011111101_011111101_011111110_011111101_011110100_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_010001110_010001110_001011101_010101010_011111110_011100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011001_011111101_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101010_011111101_010001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011100_011111101_010001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111100_011111111_011111110_001010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_011111110_011111101_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111110_011010111_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111010_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_45 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111011_010110000_001001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001001_011111110_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_010001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101100_011111110_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_011111000_011111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010101_011111110_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000101_011111110_011001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011110000_011111110_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001010_011111110_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100101_011111110_011111110_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011001111_011110101_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_011011000_011111110_010101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111110_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011111110_011111110_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111000_011111110_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011110000_011111110_011011110_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011001110_011111110_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011001011_011111110_011111110_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_011111110_011111110_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011111110_011111110_010101101_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_011111110_011111110_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_011001100_011111110_011011010_000011001_000000000_000000001_000001100_000001100_000001100_000000111_000001100_000001100_000000001_000000000_000110000_011111110_010101101_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010110_011111110_011111110_011100001_010010100_010010100_010010111_011111110_011111110_011111111_011001101_011111110_011111110_001011010_000001101_001110110_011111110_010011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101001_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011011010_011100001_011010011_011111110_011001011_011100000_011111110_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101011_011111110_011111110_011100000_011001001_010111101_010111101_001111011_001000111_001000111_000010001_000011011_000000111_001000101_010110010_011111110_011001111_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000110101_000110101_000011100_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010100_011111110_010010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_000100011_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_46 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111111_010100101_000000000_000000000_000000000_000000000_000000000_000000000_001000110_011111110_010110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000011_011111110_010011001_000000000_000000000_000000000_000000000_000000000_000000000_001101010_011111110_011111001_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011000_011111110_001101001_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111110_011110000_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011100001_011111110_001010100_000000000_000000000_000000000_000000000_000000000_001010101_011101001_011111110_011010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111010_011111110_011111110_000101110_000000000_000000000_000000000_000000000_000001000_010111010_011111110_011111110_011001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111010_011111110_011111110_000001001_000000000_000000000_000000000_000000000_010010010_011111110_011111110_011111110_001111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010110_011111110_011111110_000001001_000000000_000000000_000000000_001111111_011111011_011111110_011111110_011101111_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011001_011111110_011111110_000001001_000000000_000000000_001011100_011110110_011111110_011111110_011111110_010110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101001_011110001_011111110_000101000_000000000_000011011_011110100_011111110_011111110_011111110_011111110_010010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100001_011111110_010101001_001100100_011110100_011111110_011111110_011111110_011111110_011111100_001000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_010110000_011111101_011111110_011111110_011110101_010100111_011111110_011111110_011001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_010110001_010010010_000100011_001101110_011111110_011111110_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001110_011111110_011111110_010000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000010_011111110_011011011_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101110_011111110_011010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011111110_001111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111001_011111110_001110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001110_011111110_001110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000010_011111110_001110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011000000_001110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_47 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_001101111_010000101_001010010_000000001_000000000_000000000_000000000_000000011_001100100_010101000_011010110_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011111101_011111101_011111101_000001011_000000000_000000000_000000100_001111111_011111101_011111101_011111101_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111000_011100111_011111101_011111101_011101110_000001010_000000000_000000000_000100101_011111101_011111101_011111101_011111101_001101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110110_011111101_011111101_011111101_010010000_000000000_000000000_000000000_000100101_011111101_011111101_011111101_011111101_010000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011101001_011111101_011111101_011111101_000111010_000000000_000000000_000000000_000100101_011111101_011111101_011111101_011111101_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_011000010_011111101_011111101_011111101_011111101_000011000_000000000_000000100_001010101_011001010_011111101_011111101_011111101_011111101_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111101_011111101_011111101_011111101_011111101_001100101_001010101_011010001_011111101_011111101_011111101_011111101_011111101_010111000_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011111101_011111101_011111101_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101010_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011111101_011111101_010111011_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111110_011111101_011111101_011111101_011111101_010110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011111000_011110010_010010101_011011100_011110010_011110010_011110010_011110100_011111110_011111110_011111111_011111110_010101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000110_010111111_011111101_011111101_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010001_011111101_011111101_011111101_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011011010_011111101_011111101_011111101_010110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101010_011111101_011111101_011111101_011111101_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011111101_011111101_011111101_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111110_011111101_011111101_011111101_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111010_011111110_011111101_011111101_011111101_011100110_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_011111110_011111101_011111101_011111101_001010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_010100000_000001011_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_48 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101001_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111100_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111101_010100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111100_011011111_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111101_011111110_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111100_011111101_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111101_011111110_000110010_000110100_010000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011111100_011010101_000110011_011000001_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011000_011111101_011111110_011111101_011001011_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011000001_011111100_011111101_011010100_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000001_011111101_011111110_010000011_000110011_000110011_000110011_010000100_011010110_011111101_011111110_011111101_011111110_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011101000_011111101_011111100_011111101_011111100_011111101_011111100_011111101_011111100_011111101_011111100_011010101_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011101010_011111101_011111110_011111101_011110100_011001011_010001110_001100110_011111110_011111101_010110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_000110010_000110010_000110010_000101000_000000000_000000000_000000000_011111101_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011000_011111101_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101001_011111100_001111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111101_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101101_011111101_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_010101100_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_49 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011111101_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011000100_011111100_011110001_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010011_011100001_001100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011111100_011111100_011111101_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011111101_011111100_011000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011111100_011111100_010110010_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111101_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011111100_011111100_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_011001011_011111101_011111100_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111000_011111101_011111101_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011111101_011111111_011010111_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000101_011111100_011111100_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011111100_011111101_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000101_011111100_011111100_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000001101_001001111_011111100_011111101_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011101010_011111100_011101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011111100_011111100_010110010_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011111100_011111100_010111101_010001101_010001100_010001100_010001100_010001100_001001111_000110000_010100101_011111100_011111100_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111101_011111101_011111101_011111111_011111101_011111101_011111101_011111101_011111111_011111101_011111101_011111101_011111101_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011101001_011111100_011111100_011111101_011111100_011111100_011110010_011010110_011010111_011110011_011111100_011111100_011111100_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_011000011_011000011_000111000_000110111_000110111_000110001_000011111_000011111_000110010_011010001_011111100_011011100_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001001_011101010_011111100_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100001_011111100_011111100_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011111101_011111101_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100101_011111001_011111100_011110010_001001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011111100_011111100_011110110_001011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011101010_011111100_010011010_001100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011111100_001010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_50 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_000101111_000101111_000101111_000010000_010000001_001010101_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_010011001_011011001_011111101_011111101_011111101_011010111_011110110_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_010001110_011110100_011111100_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011010101_010101010_010101010_010101010_010101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_010000100_001001000_000000000_000111001_011101110_011100011_011101110_010101000_001111100_001000101_000010100_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_011001110_011111101_001001110_000000000_000000000_000100000_000000000_000011110_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_010110001_011111101_010000100_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_010000101_011111101_011101001_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011111101_011011111_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010110_011111101_010101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101010_011111101_011110110_001111111_000110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111101_011111101_011111101_011111011_010010011_001011011_001111001_001010101_000101010_000101010_001010101_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001011_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011101000_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_000110101_011011010_011011110_011111011_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111100_001111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_001001000_011001000_011111101_011111101_011111101_011111101_011111101_011111101_011111101_010101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111000_011111101_011111001_010011000_000110011_010100100_011111101_011111101_010101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011111101_011111101_011111101_010111100_011111100_011111101_011111101_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010100111_011111101_011111101_011111101_011111101_011111010_010101111_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_010110100_011100111_011111101_011011101_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_010010101_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_51 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_010000100_011010110_011111101_011111110_011111101_011001011_010100010_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_010001110_011001011_011001011_011111101_011111100_011111101_011111100_010010111_001000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011110100_011001011_010001110_001100110_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101100_011111100_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011011111_011101010_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111010_011111101_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011111110_001011011_000110011_000110011_000110011_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011011111_011111101_011111100_011111101_011111100_011111101_010101100_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011010110_011111101_011001011_010100010_001100110_001100110_011001011_011011111_011111110_011111101_000110011_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_011111101_010101011_000000000_000000000_000000000_000000000_000000000_000010100_001110000_011000000_011111101_011010100_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011001011_011101010_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011010101_011101000_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111110_011001011_011101010_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011010101_011111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011001_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011101001_011010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_010101101_011110100_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011111101_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000010101_001100110_001100110_010110111_011101001_011010100_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011111111_011111101_011101010_010011000_010011001_011000001_010101101_011111101_011111110_011111101_011111110_011010101_010001110_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_010010111_010010111_011101000_011111101_011010100_011000000_010010111_010000011_000110010_000110010_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_52 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_010011000_011101101_011111110_011111110_011111111_011111110_011111100_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010111_010100100_011101101_011111101_011111110_011011010_010001010_001010011_000100111_010011010_011111110_010000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001010_011110110_011111101_011111110_011011000_010100111_000110110_000000101_000000000_000000000_000000000_001100100_010111111_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101001_011111110_010101001_000110101_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000100011_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101110_011111110_001011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011110101_011011101_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001110_011111110_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010111_011111110_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011110010_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_011110000_011001011_000101100_000101100_000101100_000101100_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_011111110_011111110_011111110_011111110_011111110_011111110_011001101_001010101_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_010111000_010101001_010000101_010000101_010100010_011010100_011111110_011111110_010100110_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_000110011_010110001_011111110_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011010001_011111110_001101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011010001_011111110_011000010_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_000000000_000001010_010001001_011110100_011111110_011000110_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_001010111_001111010_010010011_011011111_011111110_011110111_001111111_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001110110_011111010_011010010_011111000_011111110_011111100_011000111_000110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001010_011111110_011111110_011111110_011111010_011001001_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_010100111_011000101_001010111_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_53 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011000001_010011000_001011100_000110011_000110011_000110011_000110011_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011011111_011111101_011111100_011111101_011111100_011111101_011111100_011111101_011000000_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111101_001100110_000000000_000010101_001100110_000111110_001100110_001100110_000111101_010110111_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101101_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_011011111_011001011_011001011_011001011_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011111110_011111101_011100000_011001011_011001011_011011111_011111110_001000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011110011_011111101_010000010_000010100_000000000_000000000_000010100_011111101_011101000_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011000_011111101_010110111_000000000_000000000_000000000_000000000_000000000_010000100_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_010010111_000010100_000000000_000000000_000000000_000000000_000000000_000110011_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_010110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000001_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_010110111_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011111110_011111101_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011011111_001100110_000000000_000000000_000000000_000000000_000000000_000010101_011001011_011111101_010000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001100_001111011_000000000_000000000_000000000_000000000_000101001_010101101_011111101_011001011_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011011111_001100110_000010101_001100110_010100011_011110011_011111101_010101011_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011101010_011111101_011111111_011111101_011111111_010101100_001010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_010000011_011000000_001101111_000110010_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_54 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_001001101_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_000111111_001110111_010101011_011110010_011110011_011001010_001100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_000010101_000000000_000011000_001110111_011001100_011111110_011111111_011100011_010000000_001101011_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_010111011_011111110_011101000_011010111_011101010_011111110_011110001_010011111_001001010_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_011011001_011111110_011111110_011111110_011111011_011011101_001101001_000100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_011000111_011111110_011111110_011111001_010100010_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111011_011111110_011111110_011000100_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_011110000_011111110_010100011_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011110_011111110_010100001_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011110010_011111000_001001100_000100010_001101011_010000110_011011010_010110001_001011101_000011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110101_011111110_011111000_011110001_011110011_011111110_011101011_011011111_011110000_011111110_011101100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_011111110_011111110_011001001_010010000_000111010_000010110_000000000_000011111_010001110_011111010_011101001_001101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_010010111_001010101_000001111_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111110_010101111_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101100_011111110_011111110_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100001_011010001_011111110_010110000_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011100100_011111110_011101001_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_001100010_010110110_011111010_011111110_011100111_001001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_000011011_000011011_001100111_001110101_010010111_011011110_011111110_011111110_011110000_010001110_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011110010_011111001_011111010_011111101_011110111_011110101_011110001_010111000_001100100_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_000110001_001000001_000100010_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_55 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_010011010_011010111_011110001_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_011101001_010110001_001000110_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110100_010010010_010010010_010010101_010110001_011100000_001110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011101_011001111_010100001_010111000_001101010_000101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_011111000_000111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_011111100_000111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_011111101_000111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011111110_000111110_000000000_000000000_000000100_000011111_000001101_000100000_000110111_000011111_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101011_011111110_000111110_000001110_001010011_011010110_011111110_011100010_011111110_011111110_011111110_010110101_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_011111110_010011010_011100001_011111011_010100111_001010100_001000110_000010111_000010111_001011011_010110011_011111010_001101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011001100_011011100_010011010_000100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011111111_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011010010_011100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011111010_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111110_011111110_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001010_011111000_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110101_011110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000001_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000001_000010010_011100101_011000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011101100_001001110_000000010_000000000_000000000_000000000_000000000_000000000_000010010_010100001_011101001_010111001_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011111110_001011010_000100000_000001100_000110111_001010101_010101000_011101010_011101010_010000001_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_010000010_011100010_011110100_011101100_011111110_011110111_010110000_001101101_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_56 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_001111011_010100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_001100111_011001010_011100001_001010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_000101000_010101011_011011111_011110000_011101100_001001010_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_001000000_010000110_011110000_011111111_011111101_010100001_000111001_000001110_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011010100_011010101_011110011_011111101_011111101_011111101_011000000_001000100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100000_011100110_011100111_011100110_010011111_001010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_001010100_001111001_000011011_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_001111110_001011110_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011001010_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011101101_011110011_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_010110100_011111111_011010010_011000001_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_000111111_000111111_010110111_010001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010101_011001100_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011100001_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_001011110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011100_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_010101101_011111110_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_001111101_011111101_011100000_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011111101_011001000_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_010000010_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_57 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_000000100_000000000_000000111_000011101_000011101_001011100_010001101_010001101_010001101_011110011_011011001_011011001_001001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_010101010_010101010_011101011_010110010_010101010_010111100_011111101_011111101_011111110_011111101_011111101_011111101_011111110_011111101_011111101_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_011101011_011111111_011111101_011111101_011111101_011111110_011111101_010111011_010101000_010101001_010101000_001010001_000111000_001001110_011111101_011100001_000101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011011111_011111101_010111111_011011000_011111101_011001011_001001110_000011100_000000110_000000000_000000000_000000000_000000000_000000000_000000100_001001110_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101010_011111110_011111111_010111111_000000000_000110011_011100010_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111101_011111101_011011000_010101010_001011111_000111001_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011111101_011111101_011111101_011111110_011111101_011111101_011100101_010000111_001000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000011100_000011100_000011100_000011100_000110101_010110010_011111101_011111110_011110111_010001010_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_001111111_011110101_011111110_011111110_010000001_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_010101100_011110111_011111110_010101100_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001010_011111110_011111101_001011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_001101000_011111101_011001110_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011111110_011111110_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011011001_011111101_011111101_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_011010010_011111110_011111101_001100011_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001100_011011111_011111101_011111110_010011000_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001001_000000100_000000000_000000000_000000000_000011010_011001101_011111110_011111110_011110010_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_010000000_000111001_001010010_010101001_011110100_011111110_011111101_011010001_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100000_011111101_011111110_011111101_011111101_011111101_011110101_010001111_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_010000000_011001100_011111101_011010111_010001100_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_58 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_001000000_011111111_010110111_011111101_010001100_001111001_001111001_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_011010100_011110000_011110000_011110000_011110110_011110110_011111101_011111100_011111100_011111100_011111100_011111100_001001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000101_011111000_011111100_011001010_011111100_011111100_011111100_011111100_011111101_011111100_011111100_011111100_011111100_011111100_011000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011111100_011111100_010100001_011101111_010101100_010101100_001100110_001101110_000100111_000100111_000100111_010100101_011111100_011110110_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011111100_011111100_001101000_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_000110101_000110101_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111100_011111100_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011110_011111100_011111100_001100000_000101001_000101001_000010011_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011010101_011111100_011111100_011111100_011111100_011001011_011001011_010100001_001101000_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_011111100_011111100_011111100_011111100_011111100_011111100_011111101_011111100_011010101_001101001_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_011111100_011111100_011111100_011111100_011111100_011111100_011111101_011111100_011111100_011111100_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_010011110_011101010_010010010_010110111_011000101_010111111_011111101_011111101_011111101_011111101_010000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_000001011_000000010_000000110_000000111_000000110_010001011_011110001_011111100_011111100_011111001_001001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011011001_011111100_011111100_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010101_011111100_011111100_011110110_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011110100_011111100_011111100_011011100_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_000001110_000000000_000000000_000100000_000110110_010111011_010111010_011110101_011111100_011111100_011111100_011010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011110_011000001_010101101_010101101_011011011_011111100_011111101_011111100_011111100_011111100_011111100_011110011_001101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011110101_011111100_011111100_011111100_011111100_011111101_011111100_011111100_011111100_011110101_001101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110001_011110001_011111100_011111100_011111100_011111101_011110110_011101110_011101110_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_010000100_011111100_011111100_001111000_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_59 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000101_010001101_011111111_011111110_011111110_011011000_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_001001000_010011010_011110100_011111101_011111101_011111101_011111101_011001011_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_001000001_010101011_011100101_011111101_011111101_011111101_011111101_011011110_001111011_001010010_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_001001000_010110000_011011101_011111101_011111101_011111101_011111101_011111101_010111100_001111010_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_010101001_011011100_011111101_011111101_011111101_011111101_011111101_010111111_010000000_000101111_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011111101_011111101_011111101_011111101_011111101_010110110_000011101_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011010111_011111101_011111101_001011110_000001011_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011111101_011111101_011111101_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_011110000_011111101_011111101_001000010_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010000_011111101_011111101_011111101_011011000_001110000_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_001011100_011101111_011111101_011111101_011111101_011110100_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100001_001011011_011001101_011111101_011111101_011110100_010010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_000100010_011010100_011111101_011110110_001011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011010110_011111101_011111100_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100100_011111101_011111101_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001000_011111101_011111101_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111101_001100000_000001100_000000000_000000000_000000111_001010101_011101000_011111101_011111101_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101011_011111101_011010011_011001001_011001001_011001110_011111101_011111101_011111101_010110010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101000_011100100_011111101_011111101_011111101_011111101_011111101_011111101_010111011_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_001110010_010000111_011000001_010111011_010000111_001101100_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_60 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011001100_011111101_010110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_010010110_011111100_011111100_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110101_011111100_010111010_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111100_001110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011110111_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011111101_011000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010110_011111101_011000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111001_001010101_001010101_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100001_011111101_001100000_000000000_000000000_000000000_000000000_000000000_010010111_011100010_011110011_011111100_011111100_011101110_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011100101_011100010_000000000_000000000_000000000_000000100_000110110_011100101_011111101_011111111_011101010_010101111_011100001_011111111_011100100_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011111100_010010110_000000000_000000000_000011010_010000000_011111100_011111100_011100011_010000110_000011100_000000000_000000000_010110010_011111100_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011111_011111100_001110001_000000000_000000000_010010110_011111101_011111100_010111010_000101011_000000000_000000000_000000000_000000000_010001101_011111100_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111001_011111100_001110001_000000000_000100110_011101101_011111101_010010111_000000110_000000000_000000000_000000000_000000000_000000000_010001101_011001010_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_011111101_001110010_000000000_010010011_011111101_010100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000101_011111100_001110001_000000000_010101100_011111100_010111100_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011111101_010101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000101_011111100_001110001_000000000_000010011_011100111_011110111_001111010_000010011_000000000_000000000_000000000_000000000_011001000_011110100_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011011110_011111100_001110001_000000000_000000000_000011001_011001011_011111100_011000001_000001101_000000000_001001100_011001000_011111001_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111001_011111101_010110011_000001010_000000000_000000000_000000000_001001100_000100011_000011101_010011010_011111101_011110100_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011010001_011111101_011000100_001010010_000111001_000111001_010000011_011000101_011111100_011111101_011010110_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_011011000_011111100_011111100_011111100_011111101_011111100_011111100_011111100_010011100_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_001100111_010001011_011110000_010001100_010001011_010001011_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_61 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_010110100_011111101_011110100_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111000_011111100_011111100_011101000_010100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011101010_011111100_010001000_000100110_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011101100_011111100_010110000_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001100_011111100_011111100_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001011_011111101_010101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011010100_011111100_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011110000_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011101_011111101_011001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100110_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100111_011111111_010110100_010001010_010110100_011111101_011111111_011111101_011011110_001100001_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100110_011111101_011111100_011111100_011111100_011111100_011010011_011111100_011111100_011111100_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100110_011111101_011110000_010110111_001011001_001000101_000000111_001000101_010101011_011111100_011111100_001010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011111101_010011001_000000000_000000000_000000000_000000000_000000000_000001101_011010111_011111100_001110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011001110_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011111100_001110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101010_011111111_011010011_000000111_000000000_000000000_000000000_000000000_000110001_011101001_011111101_001110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011111_011111100_010011010_000001001_000000000_000000000_000011110_011000101_011111100_011111100_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011100011_011111100_010011010_001000110_001010001_011100100_011111100_011100011_010000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011100011_011111100_011111100_011111101_011111100_010111001_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_010110011_011111100_010111110_001110101_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_62 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011111111_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011111111_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011111111_001110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011111111_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_011111111_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011111111_011100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111111_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000111001_001010110_001010110_010001101_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101010_011111111_001010110_000000000_000000000_000000000_000000000_000000000_000111001_011100010_011111111_011111111_011111111_011111111_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101010_011111111_001010110_000000000_000000000_000000000_000000000_000000000_010101010_011111111_011111111_001110010_000111001_011100010_011000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101010_011111111_001010110_000000000_000000000_000000000_000000000_000111001_011111111_011111111_001010110_000000000_000000000_010101010_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101010_011111111_001010110_000000000_000000000_000000000_000000000_010101010_011111111_001010110_000000000_000000000_000000000_010101010_011111111_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111111_001110010_000000000_000000000_000000000_000011101_011111111_011000110_000000000_000000000_000000000_000000000_010101010_011111111_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011111111_011111111_000000000_000000000_000000000_010101010_011111111_001110010_000000000_000000000_000000000_000000000_011000110_011100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_011111111_001110010_000000000_000000000_010101010_011111111_001010110_000000000_000000000_000000000_001010110_011111111_001110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111111_011111111_010101010_000111001_011111111_011111111_000011101_000000000_000000000_001010110_011100010_011100010_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011100010_011111111_011111111_011111111_011111111_001010110_001010110_010101010_011111111_011111111_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_010001101_011111111_011111111_011111111_011111111_011111111_011111111_011000110_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011111111_011111111_010001101_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111111_011111111_010101010_010101010_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011100010_010101010_001110010_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_63 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_010011100_011110110_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011011001_011111101_011111010_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111111_011111101_011111101_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_011110110_011111101_011000011_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011111110_011001000_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100100_011111110_011110001_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_010110111_011111101_001101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011111101_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_010000110_011011000_000100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_011110100_011111101_001001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011001_011111110_010110111_000001000_000000000_000000000_000000000_000101001_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_001001110_000000000_000010000_010001100_011010110_011110001_011011001_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_011111110_011110111_000110110_000000000_010000111_010011000_010100110_011111101_011111101_011011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000011_011111110_010110100_000000000_000000000_000000000_000000000_000001100_011011111_011111101_011111101_001001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000011_011111110_001100011_000000000_000000000_000000000_000000000_000010100_011111101_011111101_011010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000100_011111111_010001000_000000000_000000000_000000000_000000000_000010100_011111110_011111110_010000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000011_011111110_010111110_001011000_000000010_000000000_000000101_001001100_011111101_011111010_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011011111_011111101_011111101_010100110_001001111_010011100_011111101_011111101_010010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_001001000_011001010_011111101_011111101_011111101_011111110_011111101_011100001_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_000111010_011001000_011010111_011000001_001001001_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_64 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_011001110_011011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011001101_011111101_011011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011001101_011111101_011111011_010001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001000_011111101_011111101_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011010000_011111101_011101110_000100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010001_011111101_011111101_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011110001_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111101_011101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_000110010_000110010_000110010_000110010_000110010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011101011_000000000_000000000_000000000_000000000_000000000_001000100_010110100_011101100_011111101_011111101_011111101_011111101_011111101_010111011_001111110_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011101011_000000000_000000000_000000000_000000000_000001101_011000110_011111101_011111101_011001100_010111111_010010100_010000000_010110000_011110111_011111101_011011110_001111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_010001100_000000000_000000000_000000000_000000000_010010000_011111101_011111101_010101000_000001110_000000000_000000000_000000000_000000000_001101100_011010111_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011010000_000000000_000000000_000000000_000000000_010101110_011111101_011111101_000111101_000000000_000000000_000000000_000000000_000000000_000000000_001110000_011111101_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011101011_000000000_000000000_000000000_000000000_010101110_011111101_011111101_000111101_000000000_000000000_000000000_000000000_000000000_000000000_001110000_011111101_011010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_011110001_000100100_000000000_000000000_000000000_010101110_011111101_011111101_010100100_000000000_000000000_000000000_000000000_000000000_000000000_001110000_011111101_001010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100111_011111101_011111101_011101000_001010101_000000000_000000000_000011001_001111101_011100101_011110100_010110101_001000000_000000000_000000000_000000000_000000000_010011101_011111101_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_011001111_011111101_011111101_011010000_000000000_000000000_000000000_000000000_001110010_011100101_011111101_011110100_001010111_000000000_000000000_000101010_011110011_011111101_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_011111101_011111101_011111010_010010110_000100100_000000000_000000000_000000000_000110100_010010100_010110101_011110101_010111000_001101010_011100100_011111101_001011111_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000001_001011000_011001111_011111101_011111101_011110010_011010011_001110000_001110000_001110000_001110000_001110110_010101100_011111101_011111101_011001111_000011010_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010000_010000111_011010010_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011010101_010000111_001010111_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000011011_010000001_010000001_010000001_010000001_010000001_010000001_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_65 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_001100101_010010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_011111100_010101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010101_011111100_010000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_010010011_011111010_010001111_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010000_011111100_001100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_011011101_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001010_011110011_001101110_000000000_000000000_000000000_000000000_000000000_000000000_000001010_001111111_011101100_011101100_010101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010111_011000101_000000000_000000000_000000000_000000000_000000000_000000000_000111100_011101100_011111100_011111100_011111100_011111000_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011110010_010100011_000000000_000000000_000000000_000000000_000000000_000001011_011000111_011111100_010101000_001000010_011010100_011111001_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011100011_000001100_000000000_000000000_000000000_000000000_000000000_010110001_011111100_010100110_000000010_000000000_011000110_011110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011011001_000000000_000000000_000000000_000000000_000000000_000111111_011111111_011001001_000010011_000000000_000000000_010010111_011110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010001_010010101_000000000_000000000_000000000_000000000_000000000_010111011_011111101_001001101_000000000_000000000_000000000_011000110_010100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010001_010111011_000000000_000000000_000000000_000000000_000000000_011011100_011100010_000001101_000000000_000000000_000101110_011110011_010000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010001_001111001_000000000_000000000_000000000_000000000_000101001_011101101_011010011_000000000_000000000_000001100_011001110_011111100_000011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010001_011000000_000000000_000000000_000000000_000000000_001001110_011111100_001101111_000000000_000000000_001110111_011111100_010101010_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010001_011100110_000000000_000000000_000000000_000000000_001001110_011111100_001101111_000000000_001001111_011111010_011111100_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101001_011111010_010000100_000000000_000000000_000000000_001001110_011111100_010100100_000101000_011011101_011101101_000111100_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101111_011100111_010011010_000001101_000000000_001100001_011111100_011111101_011111100_011111100_001111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011100010_011111100_011000001_010111011_011101100_011111100_011111101_011111100_011111100_001010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_010001110_011110011_011111100_011011011_010001110_010011101_011011111_001100100_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_66 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_010101000_010001100_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011000110_011110011_011111110_011111110_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001011000_011111101_011111110_011111110_011111110_011111110_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011111110_011111110_011111110_011111110_011001111_010000110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_010110000_011111110_011111110_011101110_001101001_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010001_011111111_011111110_011111011_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011010110_011111110_011100001_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000111_011111110_011111011_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101011_011111111_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101011_011111110_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_011111011_011100010_000101000_000000000_000000000_000000000_000000000_000010001_001100100_011000101_010101011_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_011111011_010110101_000000000_000000000_000000000_000000000_001001011_011111001_011111110_011111110_011111110_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101011_010110101_000000000_000000000_000000000_000010011_011011101_011111110_011111110_011111110_011111110_011101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101011_010110101_000000000_000000000_000000000_001101100_011111110_011111110_011110100_010100111_011011000_011101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101011_011001100_000001010_000000000_000000010_010111010_011111110_011110010_001001001_000001010_011001101_011101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011111111_010000110_000001000_000000110_011111110_011111110_001110111_000000000_001011100_011111110_010101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100111_011111110_011111110_010101111_001001000_011111110_011111110_010010011_001101001_011111010_011111110_000011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_010110101_011111101_011111110_011111110_011111110_011111110_011111110_011111110_011111110_010110111_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011111110_011111110_011111110_011111110_011111110_011101010_010111000_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_001001000_011101110_011101001_010010110_010000101_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_67 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_010101110_011111110_001011101_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_011000111_011111101_011111101_011111101_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011111101_011001000_001100000_011001110_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100001_011100110_011111101_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011111101_011101100_001000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111101_010010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_011101110_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111101_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011111101_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011101_011111101_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_001001100_011001010_010011011_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011110_011111110_011111110_000111100_000000000_000000000_000000000_000000000_000000001_001010010_011010001_011111110_011111110_011011100_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011101_011111101_011111101_000111100_000000000_000000000_000000000_000000000_001010010_011111101_011111101_011111101_011111101_011111101_011011001_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111101_011111101_000111100_000000000_000000000_000000000_000010010_011010001_011111101_011100111_010001000_001100000_011011000_011111101_001101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111101_011111101_000111100_000000000_000000000_000000000_010010000_011111110_011010110_000100000_000000000_000000000_011000010_011111101_010011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011101001_011111101_001011001_000000000_000000000_010100101_011111010_011110110_000011111_000000000_000000000_000000000_011000010_011111101_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011111101_011101100_001001000_000011100_011101101_011111101_001110100_000000000_000000000_000001110_001100110_011101111_010111100_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100001_011100101_011111101_011101101_011100000_011111101_011111101_000000000_000000000_000110101_010101111_011111101_011111101_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011100111_011111101_011111101_011111101_011111101_011010101_010100110_011110000_011111101_011111101_010010000_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101111_011101001_011111101_011111101_011111101_011111110_011111101_011111101_011101000_001110100_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_001110100_010000100_011111000_011111110_011110010_010000100_000110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_68 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_010001101_011100000_001001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111010_011111101_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111110_010101011_001110011_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110100_011111000_011110100_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011011011_011111101_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001110111_011111110_010101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100111_011111101_011010100_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011000100_011100100_000101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010101_011111101_010101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000010_011111101_001100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011111111_010101110_000000000_000000000_000000000_000000000_000110010_001100001_000111011_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110100_011111110_010000111_000000000_000000000_000110101_011010111_011110111_011111101_011111101_010111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000011_011111110_010000111_000000000_001011000_011101011_011111110_011011000_001101011_010101100_011111101_001000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000011_011111110_010000111_001011000_011111011_011111101_010011010_000011001_000000000_010001000_011111101_010101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000011_011111110_010010110_011101011_011101101_001110110_000000000_000000000_000000000_010001000_011111101_001100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111111_011111110_011111110_010011010_000000000_000000000_000000000_000000000_010001001_011111110_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011010000_011111101_011111101_001111100_000000000_000001101_000010100_000010100_010110111_011110101_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111111_011111101_011111101_011110001_010101111_011100000_011111101_011111101_011111101_001111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001101110_011110001_011111101_011111101_011111110_011111101_011111101_011011000_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_010100011_011111101_011111110_011111101_011011110_001011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_69 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_010011101_011110001_011110111_010000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_001010111_011110001_011110001_011000110_011011110_011111101_010011000_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_010101000_011111101_011110011_000101001_000000000_000010000_010110010_011111110_001101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011111101_011001111_000100111_000000000_000000000_000000000_000110100_011101011_001111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011110011_011110000_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011010001_011110011_001000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011010001_011111101_010010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001000_011111110_011100001_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011101110_011111110_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011111101_011001010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011111110_010110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_010000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011111101_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011101110_011111101_010000001_000000000_000000000_000000000_000000000_000001100_000010011_000010011_000010011_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011101110_011111101_010110101_000000000_000000000_000101000_001111100_011100100_011111101_011111101_011111101_011100011_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001101_011111110_011001010_000000101_010011001_011111110_011111110_011111111_010111010_010111111_011111110_011111110_011001010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011010_011111101_011111110_011101101_011111010_011011111_001101100_000010010_000000010_000000011_011001011_011111101_011111110_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_010010001_011111110_011111101_011111101_001111101_000000000_000000000_000001000_000110010_011100010_011111101_010010010_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011010000_011111101_011111101_011111001_011000111_011001000_011010011_011111101_011111011_010101001_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_001111100_010101111_011111101_011111101_011111110_011111101_011001111_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_70 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_010111001_010011111_010010111_000111100_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011110_011111110_011111110_011111110_011111110_011110001_011000110_011000110_011000110_011000110_011000110_011000110_011000110_011000110_010101010_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_001110010_001001000_001110010_010100011_011100011_011111110_011100001_011111110_011111110_011111110_011111010_011100101_011111110_011111110_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_001000010_000001110_001000011_001000011_001000011_000111011_000010101_011101100_011111110_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010011_011111101_011010001_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011101001_011111111_001010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000001_011111110_011101110_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111011_011111001_011111110_000111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000101_011111110_010111011_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_011001101_011111000_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111110_011111110_010110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_011111011_011110000_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011011101_011111110_010100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_011001011_011111110_011011011_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011111110_011111110_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011100000_011111110_001110011_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000101_011111110_011111110_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_011110010_011111110_011111110_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111110_011111110_011011011_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_011111110_011001111_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_71 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001010_011111001_011111110_011111110_011111110_011110101_010100111_010100111_010001000_000011001_001010000_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101000_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111001_011111110_011111100_011000101_001110001_001000111_000100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001100011_010000111_001101001_001101001_001110010_011000000_011000000_011000000_011101001_011111110_011111110_011111110_011111110_011111110_011110110_010000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_001110010_001110010_011001011_011111110_011111110_011111110_011110000_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_000100011_010011011_011111110_011111110_010000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011111110_011110001_000100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110011_011111110_011111110_001110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011110011_011111110_011110000_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101111_011111110_011111110_010001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011110011_011111110_011110100_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_010110000_011111110_011111110_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111110_011111110_011011100_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111101_011111110_011110011_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111111_011110001_011111110_011111110_001010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_011110011_011111110_011111110_010010011_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_001101111_011111110_011111110_011001011_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111010_011111110_011111110_011111110_001010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011101101_011111110_011111111_011000010_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011111110_011111110_011000010_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100111_011100110_011000001_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_72 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_000000000_000000000_000000000_000001011_001011100_010101101_011111101_011111110_011111101_011111110_011111101_000111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001110_000000000_000010101_001100110_011010101_011111100_011101001_010010111_010000011_010000011_011111101_011111100_010001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_010011000_010011000_011010110_011101001_010110111_001100110_000000000_000000000_000000000_000000000_010000100_011111101_011111111_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011110011_011111101_011111100_010000011_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011010100_011111101_010000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011001011_001100110_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011111111_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111101_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111110_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111101_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100011_011111110_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011111101_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011011111_001111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101001_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011111101_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011111110_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011011111_011101001_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111101_010110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011111100_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_73 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100100_011010011_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000110011_001111001_001111001_011100010_011111101_011101000_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_011101011_011111001_011110000_011110000_011110000_011110000_011110000_011110001_011110101_011111100_011111100_011111100_011111100_011111100_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_010110111_011111100_011111100_011111100_011111100_011111100_011111101_011111100_011111100_011111100_011111100_011111100_011111100_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_000100111_000100111_000110101_001011111_000100111_000100111_000100111_000100111_011011011_011111100_011111100_011000101_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_011110100_011111100_011010001_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111010_011111100_011111100_011000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011110100_011111100_011111100_010110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011110001_011111100_011111100_001111110_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011000101_011111100_011111100_011111000_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011000100_011111101_011111100_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011000101_011111101_011111111_011111101_010011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_001111011_011111100_011111100_011111101_011111100_001100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011010_011111100_011111100_011111100_011111101_000100101_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011000110_011111100_011111100_011010001_001101110_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_010110000_011111100_011111100_011111000_001011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_001101011_011111100_011111100_011111100_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101011_011111100_011111100_011111100_011101001_000100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011011001_011111100_011111100_011111100_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011001_011111010_011111100_011111100_011011101_000100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010101_011011001_011011001_001001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_74 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_010011100_010010100_001011001_001010001_010011100_011111111_011111110_011111110_011111110_011011000_010011100_010010100_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011001111_011111110_011111101_011111101_011111101_011110101_011101010_011000011_011101001_011101001_011101001_011110110_011111101_011110001_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100110_011111101_011111110_011111101_011111101_010000000_000110000_000000000_000000000_000000000_000000000_000000000_000110000_011100010_011111101_001010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_010101110_011111011_011111101_011110100_001111100_000010011_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010110_011111101_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011111101_011111101_010110001_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_011110100_011111101_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011000011_001011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110011_011111110_010011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011111110_011111011_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_011111110_010100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100101_011111000_011111110_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001101_011111101_010101011_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011101111_011111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_001011100_011111101_011111101_011010111_011010110_011010110_010110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_010100111_011111101_011111101_011111101_011111110_011111101_011111101_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001001_011111101_011111101_011111101_010111001_001110101_000100010_000010011_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110111_001001001_011000001_011101101_000100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010000_011111110_011010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111101_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111101_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011000001_000100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_75 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_001100001_010110101_011111110_011111111_011011101_001101010_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_010000000_011010101_011110101_011111110_011111110_011110110_011101111_011111110_011111110_001011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_010010111_011101111_011111110_011111110_011011110_011001100_010111101_001000110_000011011_011010111_011111110_001100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011111000_011111110_011101001_000101000_000001111_000000000_000000000_000000000_000000000_001100000_011111110_001101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111001_001001000_000100001_000000000_000000000_000000000_000000000_000000000_000000000_001001100_011111110_010111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011110_011111110_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111100_011111110_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_011001011_010101110_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111110_001111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_011011111_011001101_011111110_001110011_000100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_011111000_011111110_011111110_011111110_011110010_010111111_001000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111110_011111110_011111000_011010001_011111110_011010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_010111010_011010000_001000111_000110001_001001010_010111111_010000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011111110_001110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_011000101_010101000_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011100001_000101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110011_011101001_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100001_011100011_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100100_001111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101000_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_76 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_010111111_011111111_010000000_010000000_010000000_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_010000000_010000000_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_010111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_001000000_010000000_010000000_010000000_010000000_011111111_011111111_011111111_011111111_011111111_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_010111111_011111111_011111111_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_011111111_011111111_010000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111111_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111111_011111111_011111111_011111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_011111111_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_010111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111111_011111111_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_77 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_011000101_011111111_011110010_010010001_011101100_011010100_010101001_010000010_010000010_010000010_001011111_001101011_010000010_001010101_001110100_001000110_001001100_000000111_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111101_011111000_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111100_001101111_001101111_001101111_001101111_001101111_001101111_010001010_011101011_011101011_011101011_011110001_011101110_011110001_011111101_011111101_011111101_011111101_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_000010010_000110000_011101111_011111101_011110010_010101010_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011111101_011111101_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001010_011110000_011111101_011011011_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101111_001010110_000101100_000101100_000101100_000001011_000000000_001001011_011101111_011111101_011101100_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010110_011100000_011111101_011111101_011111101_011111101_011000001_010101110_011101110_011111101_011111101_010101101_000110010_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_011001110_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011011101_010110100_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_001000100_010000000_010011011_011101101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_011111101_001100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011101101_011111101_011111101_011000110_010001110_000111101_000111101_000111101_000111101_000111101_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_010101111_011111101_011111101_010011110_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010110_011111101_011111101_001100010_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011110000_011111101_010011111_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100001_011110001_011111101_011001101_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010111_011111101_011101010_000111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_011110101_011111101_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011110111_011111101_011101010_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_011111001_011111101_011101100_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011111101_011111101_010011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_78 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_000001101_000001101_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011110_011111011_011111011_011111011_011100101_011110100_011111011_011111011_011111100_011001111_011010000_011110001_011101010_010110111_010000000_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110101_011111101_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111001_010110111_010100000_001100100_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_000001101_000001101_000001101_000001101_000001101_000001101_001011000_001100011_010001101_001110011_010001010_011101111_011111110_011111110_011111110_011111110_011111111_001101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_000110110_010101000_011101101_011111110_011111110_011111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011101101_011111110_011111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011011111_011111110_010110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011111111_011111110_001101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101010_011011110_011111110_010011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011011111_011111110_011101110_001000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011010010_011111110_011111101_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_010111111_011111110_011111100_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001011_011111110_011111110_010111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_011110011_011111110_010111110_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011100100_011111110_011100101_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011010000_011111110_011111110_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_011000011_011111110_011111110_010000111_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011111110_011111110_010100101_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000001_011111110_010110010_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_001000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_79 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011100010_011010110_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_000011001_000011001_000010011_000000000_000000000_000000000_000001011_000011001_000001101_000011001_000011001_000110000_011011111_011111101_011110101_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010001_011111101_011111101_011100110_001000001_010000111_010011101_011000111_011111101_011010001_011111101_011111101_011111101_011111101_011111101_010010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011010100_011011101_011001101_011011011_011100110_011111101_011111101_011111101_011111110_011111101_011111101_011111101_011111101_010110101_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_000011000_000000000_000010101_000100110_001001000_001001000_001001000_001001000_001001000_010111000_011111101_011101111_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_010111001_011111101_001100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111100_011111101_011111101_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010001_011111101_011101011_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_001101110_001101110_001101110_011000000_011111101_011111001_010001111_001101110_001101110_010100111_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011111100_011111101_011111101_011111110_011111101_011111101_011111101_011111101_011111101_011111101_011111101_001010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101001_011100111_011110010_011110100_011111110_011111110_011110110_010111000_010010101_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011111101_011111010_001001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011111101_011011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011110_011111101_011011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000101_011111101_011011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100010_011111101_010110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_001100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_001100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_001100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010001_011110010_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_80 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_000101111_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_001101100_011111001_011111101_011111101_011010000_011001111_011001111_011001111_010010101_001000001_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010111000_011111110_011111101_011111101_011111101_011111110_011111101_011111101_011111101_011111110_011111101_011010101_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011001011_011111110_011111110_011000111_001111111_001111111_000111100_001011101_001010100_001000100_010010111_011011110_011111110_010100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001010_011111101_011111101_011000111_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011111101_011010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001010_011111101_011111101_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001010_011110001_011111101_011010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101001_011111101_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011100101_011111101_011111101_010100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010101_011111110_011100101_000101000_000000000_000000000_000000000_000100110_010011001_011111110_011111110_011111110_010110100_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011000110_011111110_011001111_000001001_000100010_001001000_011101011_011111101_011111101_011100000_010001011_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011010011_011111101_011010111_011110000_011111110_011111101_011101010_010000000_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011100101_011111101_011111101_011111101_011100100_001001101_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_010101010_011111110_011111110_011111110_011111110_011111110_011111110_001110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_010000010_011100110_011111110_011111101_011111101_010111001_001110011_001000000_011010011_011111101_011111000_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100110_011101000_011111101_011111101_011110111_010100010_000101110_000001101_000000111_001011011_011110101_011111101_011111110_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111101_011111101_011111101_011010010_001011101_001111111_010011111_011001100_011111101_011111101_011111101_011100100_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011110001_011111110_011111111_011111110_011111110_011111110_011111110_011111110_011111110_011100100_000100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_001110011_010001100_011001110_011001110_011001110_011001111_011001110_001111011_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_81 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_001001011_000000000_001100010_010111001_010110010_001011110_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_001101111_011000011_011101110_001011110_000000000_011010000_011111001_011111110_011111110_001110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_000110010_001101011_011000101_011110110_010110111_000011001_000000000_000000000_001010001_011110101_011111110_011111001_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_001010100_011100110_011111110_011111110_011011101_001010110_000000000_000000000_000000001_001111101_011111101_011111110_010110010_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000101_011111110_011111110_011011001_001110110_000000100_000000000_000000000_000111110_011001010_011111110_011110001_010000011_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101011_011110100_011111110_011010101_000101101_000000000_000000000_000000000_000111110_011110000_011111110_011011100_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011110110_011111110_011010001_000110001_000000000_000000000_000000000_000011111_011110001_011111110_011011101_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011111110_011111110_000110111_000000000_000000000_000000000_000010001_011000110_011111110_011011010_000011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011011011_011111110_011101001_010010000_000100111_000101010_011001100_011111110_011001101_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110011_011111000_011111110_011111110_011110100_011101001_011111110_011011111_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_001010100_010101000_011110101_011111110_011111110_011111110_011001111_001110011_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011101100_011111110_011100110_010100011_011101101_011110100_011010011_001010000_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111110_011111110_001100011_000000000_000000000_000100101_011100001_011111110_010000010_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_011111110_011100101_000001100_000000000_000000000_000000000_000000010_010101010_011111110_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100000_011111110_011111110_000010010_000000000_000000000_000000000_000000000_001010001_011111110_011000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010000_011111110_011111110_000010010_000000000_000000000_000000000_000000000_010000011_011111110_001110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_011010110_011111110_001001110_000000000_000000000_000000000_000000001_010110111_011110100_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011111101_011011111_000011000_000000000_000000010_001111110_011111110_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010111_011101110_011011110_001110111_010110001_011111110_011011001_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_010011010_011000100_011000100_001100101_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_82 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_001111111_011010001_010110010_010000110_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_010110010_011110111_011111101_011111101_011111101_011111110_010100111_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111010_011101011_011111110_011011000_001101011_001001110_001110011_011111110_011111101_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011101101_011111101_010000011_000001010_000000000_000000000_000110101_011111110_011111101_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_010110111_011111101_010001011_000000000_000000000_000000000_000011111_011011001_011111110_011001000_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011001110_011111110_000111010_000000000_000000000_001100110_011111110_011111110_011011010_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101111_011111101_001000010_000100011_001111101_011110001_011111101_011001000_000111001_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101111_011111101_011011111_011100000_011111101_011111101_011111101_011000001_010010010_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001010_011111101_011111101_011111110_011110101_010111001_011100111_010001010_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_011110101_011111101_011111110_011111101_011000000_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_010100100_011111110_011111111_011101110_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101100_011110001_011111101_011001111_011001001_011111101_011100010_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011110001_011111101_011000011_000110000_000101001_011110001_011111101_010010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_010011000_011111110_011111010_001110100_000001001_000000000_000000000_001001000_011111101_011111010_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_011111101_011111110_001111001_000000000_000000000_000000000_000000000_000010100_011111101_011111101_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000101_011111110_011011010_000001111_000000000_000000000_000000000_000000000_000101011_011111110_011110100_000101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000011_011111010_011111101_001000100_000000000_000000000_000000000_000001000_001100111_011101000_011111101_001111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011111101_011111101_001001111_000010010_001001111_010101000_011001101_011111110_011111101_010101000_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_011100011_011111101_011111110_011101110_011111101_011111101_011111101_011000000_001101101_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101111_011100110_011111110_011111101_011011110_001100111_000111010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_83 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_001111001_001111001_001111001_010111110_011111111_011111101_011111101_011111101_011111101_011111101_011101000_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000100_011110000_011110010_011111100_011111100_011111100_011111100_011111101_011111100_011111100_011111100_011111100_011111100_011111100_001011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011111000_011111100_011111100_011111100_011111100_011111100_011111100_010011111_010011110_011000001_011111100_011111100_011111100_011011000_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011110000_011111100_011111100_010110000_000100111_000100111_000100111_000000000_000000000_000001111_001101011_011111100_011111100_010110110_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010101_011111100_011111100_011000011_000011001_000000000_000000000_000000000_000000000_001101110_011011000_011111100_010101110_000011001_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111000_011010101_011111100_011111100_011000100_000110011_000000000_000011010_010110100_011110101_011111100_011101110_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101101_011111100_011111100_011111100_011111000_010101101_011010011_011111100_011111100_011101111_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_011000100_011111100_011111100_011111100_011111100_011111101_011111100_011110010_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_001111111_011110111_011111100_011111100_011111101_011111100_010100011_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011010_011111100_011111100_011111101_011111100_011111100_001101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011001100_011111101_011111101_011111111_011111101_011111101_010101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100001_011111100_011111100_011000011_010010010_011110111_011111100_011001110_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_011110100_011111100_011110000_000001100_000000000_001010001_011110010_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100110_011111100_011111100_001111110_000000000_000000000_000000000_011100010_011111100_011110010_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_011101110_011111100_011111100_001101010_000000000_000000000_000000000_001111010_011111100_011111100_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_011101110_011111100_011111100_001101010_000000000_000000000_000000000_001011110_011111100_011111100_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111010_011111100_011111100_001111111_000000000_000000000_000100111_010111101_011111100_011110001_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100111_011111100_011111100_011110111_010100000_010100001_011110111_011111100_011111100_010101011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010111_011000101_011110111_011111100_011111100_011111101_011111100_011110111_011000100_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001100_001111110_011111100_011111101_001111110_001001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_84 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_010101011_011111111_011111110_011111111_010111001_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_000111111_000101101_000000000_001110111_011110111_011111001_010111111_010111111_011100110_011111110_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010111_011101110_011111110_011110110_011100100_011110010_001111000_000011001_000000000_000000000_001001101_011111110_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001001_011111110_011111110_011111110_011111110_011000100_000000000_000000000_000000000_000000000_001111100_011111110_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111011_011111110_011111110_011110111_010110011_001000100_000000000_000000000_000000000_000101100_011111001_011111001_000100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_010101010_011111110_011101011_000110011_000000000_000000000_000000000_000101010_011101000_011111110_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011100011_011111110_011101011_010001111_000000000_000101011_011100111_011111110_010110010_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011110_011111101_011111110_010110001_001000111_011100111_011111100_010011010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111110_011111011_011111011_011111110_010110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101111_011111000_011111110_011111110_010111111_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110100_011011101_011111110_011111110_011111110_010111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110100_011101100_011111001_010111000_011001011_011111110_011101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_011101011_011111100_001010101_000000000_001000110_011111110_011111001_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001100_011111110_010001100_000000000_000000000_000101101_011111110_011111110_010000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011111100_011111000_000011111_000000000_000000000_000010010_011100011_011111110_011010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111110_011000010_000000000_000000000_000000000_000000000_010000000_011111110_011111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_011111110_010101001_000000000_000000000_000000000_000000000_010000110_011111110_011111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011010011_011111100_001110011_000011011_000110000_010000100_011110101_011111110_011000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111110_011111110_011111110_011111110_011111110_011111110_011100111_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_001101110_011000010_011111110_011111110_011111110_010101001_000010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_85 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_010001001_011011000_011111111_011110101_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_001001100_011010100_011111101_011111101_011111101_011111101_001010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100111_011010100_011111101_011111101_011111101_011111101_011111011_011111101_010000100_000000000_000001111_010001101_011011110_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011100100_011111101_011111101_011101111_010011101_001100110_000111011_010100001_001010110_000111011_011001110_011111101_011111101_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_010011101_011111101_011111010_010101100_001000100_000000000_000000000_000000000_000000110_001100110_011010110_011111101_011111101_010111010_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011001_011111101_011111010_001011110_000000000_000000000_000000000_000000000_000000100_001111011_011110101_011111101_011101100_001101011_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011110_011111101_010101100_000000000_000000000_000000000_000000000_000100010_011000000_011111101_011111101_011101011_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011110_011111101_001011010_000000000_000000000_000000000_000101011_010101000_011111101_011111101_011000100_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011110_011111101_010101000_000001001_000000000_000000110_010110011_011111101_011111101_011110101_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000111_011111101_011111101_011001110_000110111_010101000_011111101_011111101_011101010_000110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011111101_011111101_011111101_011111101_011111101_011111101_010101011_000100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000001_001010001_011001100_011111011_011111101_011111101_011111101_001100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011110101_011111101_011111101_011111101_011010100_000100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011111101_011000001_010111101_011111101_011111101_011101100_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011011011_011110011_000000100_000000100_010100100_011111101_011111101_001001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101100_011111101_011110011_000000000_000000000_000000110_001110110_011111101_011001011_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011010_011100011_011110111_000101000_000000000_000000000_001100011_011111101_011101011_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000001_011111101_011111011_011111001_011001011_011111100_011111101_011011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_010101111_011111101_011111101_011111101_011111101_011111101_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_010010001_011100100_011111101_011100110_000111100_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_86 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011010110_011111101_011111110_011010101_010000100_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_010100010_011111101_011111100_011111101_011111100_011111101_010101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011111101_011111110_010000011_000111110_001100110_011000001_011111101_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101001_011111100_010101100_000001010_000000000_000000000_001000111_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111110_011111101_000000000_000000000_000000000_000000000_000110011_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001110_011111101_010101011_000000000_000000000_000000000_000000000_001011100_011111100_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001011_011111110_001011011_000000000_000000000_000000000_000101001_011010110_011111101_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011110011_011101001_000011110_000000000_000000000_000101001_011110011_011111101_011010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011111101_011101010_000011110_000000000_000000000_010101101_011111101_011111110_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_011111100_011111101_010101100_000010101_010110111_011111101_011111100_011111101_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110111_011111110_011111101_011111110_011111101_011111110_010101100_011111110_011111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111101_011010101_011111100_011111101_011111100_010000011_000001010_010000011_011111100_001111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011111101_011111110_000110010_000000000_000000000_000110011_011111101_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011101001_011111100_010101100_000001010_000000000_000000000_000110011_011111100_011011111_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_000000000_000000000_000000000_000000000_000110011_011111101_011001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011111101_011111100_000000000_000000000_000000000_000000000_001011100_011111100_010100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100111_011111111_011111101_000000000_000000000_000001011_010101101_011111111_011101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100110_011111101_011111100_000101001_000101001_010101101_011111100_011010101_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011101010_011111101_011111111_011111101_011111111_010101100_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000111_011111100_011111101_011010100_001011011_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_87 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001001_000111000_001001111_011110000_010100001_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_000001010_000110000_011000011_011111110_011111110_011111110_011111110_001110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110100_001011011_011111010_011111110_011111110_011111110_011111110_011100001_011101001_011110110_001001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_001110111_011110111_011101000_011111110_011111110_011101011_010010111_000100011_000010100_010110001_011111110_010101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001111_011100111_011111110_011111110_011111110_010011111_000000010_000000000_000000000_000010000_011111110_011110111_001010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011001110_011111110_011111110_011111110_010100001_000000001_000000000_000000000_000100001_011011101_011100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110101_011010101_011111110_011111110_011111110_000000101_000000000_001110101_011110100_011111110_010100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111011_011011000_011111110_011111110_010110101_000011100_010101111_011111110_010111100_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001101_010101110_011111110_011111110_011010000_011111110_011111110_001101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_010001101_011111110_011111110_011111110_010110100_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_011111011_011111110_011111110_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011010001_011111110_011111110_011111110_011110011_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_010000011_011111110_011111110_011110000_011001110_011111110_010101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010000100_011111110_011111110_011110001_000100100_000010100_011001001_011100111_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_010101010_011111110_011111110_011111110_001000011_000000000_000000000_001101010_011111110_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001100_011111110_011111110_011110010_001100010_000000010_000000000_000000000_000000101_011000011_011101101_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110011_011111110_011111110_011011100_000100100_000000001_000000000_000000000_000000000_001001110_011111110_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010011_011101100_011111110_011111110_011111110_010111111_010111110_010111110_010111110_011010000_011111110_010101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101101_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_010101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011100011_010011010_001000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_88 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_000100010_001110100_010001111_011001110_011111101_011111101_010111010_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001010_011110110_011111100_011111100_011111100_011111101_011111100_011111100_011111100_010100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_011110011_011111100_011111100_011111100_011111100_011110000_010011001_010011001_010100010_011000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100001_011111100_011111100_011101111_010010100_000011000_000001001_000000000_000000000_000000001_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_011111100_011110101_000100010_000000000_000000000_000000000_000000000_000000000_000000000_000001101_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_011111100_011111010_001110100_000000000_000000000_000000000_000000000_000000000_000111000_011010010_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101111_011110101_011111100_011111001_001110101_000000010_000000000_000001000_010010010_011110010_011111010_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011001001_011111100_011111100_001110111_000111011_011011111_011111100_011111100_010110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_010111101_011111100_011111100_011111101_011111100_011111100_010011010_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011001_011100000_011111100_011111101_011111100_011010001_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010100_011010010_011111101_011111101_011111111_011111101_011010010_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111110_011110110_011111100_011111100_011111100_010001011_011101000_011111100_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011001_011111100_011111100_011111100_010100001_000000000_000011111_011011001_011101111_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010010_011111100_011111100_011010100_000010100_000000000_000000000_001100000_011111011_011000110_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_011111100_011111100_001101000_000000000_000000000_000000000_000000000_011011010_011111100_000110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000110_011111100_011101101_000101011_000000000_000000000_000000000_000000000_010101011_011111100_010001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111100_011100101_000100101_000001010_000001100_000001100_010010010_011111011_011111100_010011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011101111_011111100_011011110_011110000_011111101_011111100_011111100_011111100_011011011_000010110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010101_011111100_011111100_011111100_011111101_011111100_011111100_011010100_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_000110100_010110000_011111100_011111101_011011111_010001110_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_89 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_001100000_001100000_001100000_010011011_011111101_010101101_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_010011010_011011100_010110100_010100001_010100001_010110101_011101100_011101100_001011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_001101110_000000000_000000000_000000000_000000000_000000000_001111111_011111011_011111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_011100001_011111011_000101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010000_011110000_011111011_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111101_011000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_010000011_010111111_010111110_010111110_000110011_000001100_000001100_000110100_011011101_011111011_001011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_001111110_001111110_011011100_011111011_011111011_010101101_010101110_011111011_011111011_011011011_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_010111100_011001100_011111011_011111101_011111011_011111011_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111011_011111101_011111011_011111011_010000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011111101_011111101_011111101_010011111_010101010_011111101_011111101_001011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011100_011000101_011111011_010111000_000111110_000000000_000001000_010011101_011111011_001011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111011_010111100_000001111_000000000_000000000_000000000_001111111_011111011_010101101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001011_011111101_011011111_000001111_000000000_000000000_000000000_000000000_001111111_011111011_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011110_011111101_001111001_000000000_000000000_000000000_000000000_000010100_011001101_011111011_001011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011000010_011111111_000111111_000000000_000000000_000000000_000100100_001110011_011111101_011100101_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_010110101_011111101_001010010_000000000_000010100_000010100_011010110_011111011_011101011_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011110_011111101_011101100_001111111_011001101_011001101_011111101_011111011_001111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110111_011111101_011111011_011111011_011111011_011111011_011100101_001000101_000001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_001011110_010101101_011010011_001011110_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_90 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_010010101_011000001_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_011100000_011111101_011111101_000010011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011101011_011111110_011111101_011111101_010100110_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010000_011111101_011111110_011111101_011111101_011111101_011101110_001110011_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_011110001_011111101_011010000_010111001_011111101_011111101_011111101_011100111_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001111_011111110_011000001_000000000_000001000_001100010_011011011_011111110_011111111_011001001_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111101_001010000_000000000_000000000_000000000_010110110_011111101_011111110_010111111_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101111_011111101_010011011_000000000_000000000_000000000_011101010_011111101_011111110_010000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111101_011010000_000101000_001010101_010100110_011111011_011101101_011111110_011101100_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_011101110_011111101_011111110_011111101_011111101_010111001_000100100_011011000_011111101_010011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_011110000_011111111_011111110_010010001_000001000_000000000_010000110_011111110_011011111_000100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_010011110_010001110_000001100_000000000_000000000_000001001_010101111_011111101_010100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111101_011100010_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_010100110_011111101_001111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110000_011110101_011111101_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110011_011111110_010101100_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_011011010_011111110_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_011111110_010100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111010_011110100_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011011111_001001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_91 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100100_000111000_010001001_011001001_011000111_001011111_000100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_010011000_011101010_011111110_011111110_011111110_011111110_011111110_011111010_011010011_010010111_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_010011001_011110000_011111110_011111110_011100011_010100110_010000101_011111011_011001000_011111110_011100101_011100001_001101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011001_011101010_011111110_011111110_010111011_010001110_000001000_000000000_000000000_010111111_000101000_011000110_011110110_011011111_011111101_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_001111110_011111101_011111110_011101001_010000000_000001011_000000000_000000000_000000000_000000000_011010010_000101011_001000110_011111110_011111110_011111110_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011110011_011111110_011100100_000110110_000000000_000000000_000000000_000000000_000000011_000100000_001110100_011100001_011110010_011111110_011111111_010100010_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001011_011110000_011111110_011011111_001101101_010001010_010110010_010110010_010101001_011010010_011111011_011100111_011111110_011111110_011111110_011101000_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010101111_011110100_011111101_011111111_011111110_011111110_011111011_011111110_011111110_011111110_011111110_011111110_011111100_010101011_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_010001000_011000011_010110000_010010010_010011001_011001000_011111110_011111110_011111110_011111110_010010110_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100010_011111110_011111110_011110001_001100011_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111010_011111110_011111110_001011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100100_011110010_011111110_011111110_011010011_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011110001_011111110_011111110_011110010_000111011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000011_011111110_011111110_011110100_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001101_011111001_011111110_011111110_010011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001100_011100100_011111110_011111110_011010000_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011111111_011111110_011111110_001000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010001_011111110_011111110_010001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011100011_011111111_011101001_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011111111_001101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_92 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_010110100_011111101_011111111_011111101_010101001_000100100_000001011_001001100_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_001000100_011100100_011111100_011111100_011111101_011111100_011111100_010100000_010111101_011111101_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110111_011111100_011111100_011100011_001001111_001000101_001000101_001100100_001011010_011101100_011110111_001000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011101001_011111100_010111001_000110010_000000000_000000000_000000000_000011010_011001011_011111100_010000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101000_011111101_010110010_000100101_000000000_000000000_000000000_000000000_001000110_011111100_011111100_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011111101_011110010_000101010_000000000_000000000_000000000_000000000_000000101_010111111_011111101_010111110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001111_011111100_011100110_000000000_000000000_000000000_000000000_000000101_010001000_011111100_011111100_001000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001111_011111100_011100110_000000000_000000000_000000000_000100000_010001010_011111100_011111100_011100011_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_011111100_011111001_011001111_011001111_011001111_011100100_011111101_011111100_011111100_010100000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001001_010110011_011111101_011111100_011111100_011111100_011111100_001001011_010101001_011111100_000111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_001110100_001110100_001001010_000000000_010010101_011111101_011010111_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111101_011111100_010100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100000_011111101_011110000_000110010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011101_011111101_010100100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011110000_011111101_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_011111101_011111100_001010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110010_011111100_011010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011001111_011111100_001110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100101_011111100_001110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011101_011001000_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_93 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_010010010_011100101_011111111_011001101_001111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_011000110_011111100_011111101_011100001_011011000_011101011_011111100_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010100_011001101_011111101_011011111_001000110_000001111_000000000_000011101_011001110_010101110_000000010_001010111_000100110_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001001_011111101_011100011_000000110_000000000_000000000_000000000_000000000_000100011_000011100_001001100_011111101_011111101_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011111011_011101011_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000101010_011101110_011111101_010101110_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000110_011111101_011000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_011101110_011111101_010100001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101001_011111101_001001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010101_011110111_011111101_001001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011111010_011111101_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000110_011011011_011111101_011110001_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001010_011111101_011111101_000101111_000000000_000000000_000000000_000000000_000000000_000000101_001001000_011111101_011111101_010001111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_011011101_011111101_001110101_000000000_000000000_000000000_000000000_000011001_001110110_011111101_011111101_011111101_000101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011110010_011111110_010111011_001101000_010010010_010011111_011011100_011110100_011101111_011111110_011100000_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001110_011001001_011111101_011111101_011111000_011010111_010011100_001000011_011110111_011111101_010011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_000111000_000111000_000110010_000000000_000000000_000100110_011111101_011111101_001001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011111101_011111101_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010101_011111101_011111101_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011110_011101110_011111101_010111111_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011111101_011111101_001110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010111_011111101_011110100_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101010_011111101_011000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011111110_011111101_010010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_94 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011111_010001100_011000001_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_010010010_011110000_011111110_011111110_011100100_000110000_001001101_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_000101011_011100110_011111110_011111110_011111110_011111110_011111110_011110001_011111110_011000101_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010101_010000010_011111110_011111110_011111110_011101111_011111100_011111110_011111110_011111110_011111110_011101101_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011010_011111110_011111110_011111001_001101000_001000111_011000110_011111110_011111110_011111110_011101010_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_010101101_011111100_011111100_011001110_000110011_001111000_011010111_011111110_011111110_011111110_011111110_010111000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110000_011111110_011111110_011010111_001010111_011110111_011111110_011111110_011111110_011111110_011111110_011011001_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000101_011100111_011111110_011111110_011111110_011111110_011111110_011101100_010000000_011000100_011111110_011111110_001110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_011000101_011111110_011111110_011110101_011101110_010000011_000010001_000101110_011110111_011111110_011000111_000001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_001011100_001011000_000101000_000000000_000000000_000001100_010101101_011111110_011110010_000100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011111110_011111110_010011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010010_011010010_011111110_011100001_000000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000101_011111110_011111110_001100011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011110010_011111110_010110011_000000011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_011011111_011111110_011100001_000011110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001101_011111110_011111111_001111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011101110_011111110_011111000_000110101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_010110111_011111110_011111110_011100111_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110001_011111110_011111110_011100110_000110000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011101111_001111110_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_95 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011011_001001001_010011101_010100011_011000011_010100011_000011011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111100_010111000_011110010_011111110_011111101_011111101_011111101_011111101_010011110_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110010_010110011_011111000_011111101_011111101_011011001_011000101_001111111_010100101_011110010_011111110_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_001110100_011101010_011111101_011111010_010100011_001010000_000000000_000000000_000000000_000000000_010110101_011111110_001101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110100_011111101_011111110_011010110_000111110_000000000_000000000_000000000_000000000_000000000_000000000_010110101_011111110_010100000_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011111110_011111110_010110110_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011100100_011111111_011111110_001111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111101_011001001_000000111_000000000_000000000_000000000_000000000_000000000_000100000_000110111_010101100_011111101_011111110_011111101_000101010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000000_011111101_011001111_001000101_000100101_000100000_000010000_001100110_010111010_011101110_011111101_011111101_011111101_011111110_010100000_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011111001_011111101_011111110_011111101_011110101_011011110_011111101_011111110_011111101_011111101_011111101_011111101_011111110_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100000_011100011_011111110_011111101_011111101_011111101_011011100_010001000_001001000_001101001_011010110_011111101_011100100_000001100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111011_001011011_000101110_000000000_000000000_000000000_000000000_000111111_011111110_011111110_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110011_011111101_011001001_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011100_011101011_011111101_001010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111111_011111101_011101110_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010010001_011111101_011001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101111_011110001_011111110_010010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110110_011111101_011110101_001010001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101110_011111110_011111101_010001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011011_011111110_011011111_001001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000111011_011000011_001000110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_96 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001110_011111110_011001100_010101100_011000111_010001100_001011011_000011011_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000100_011011110_001010001_001001010_010011001_010111001_011101101_011101101_011111010_011000010_000011101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100110_011000100_000000000_000000000_000000000_000000000_000000000_000000000_001110011_001010001_000001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010101_010011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000111_011011100_001110011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100010_011110110_010000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010101000_011110110_000010101_000000000_000000000_000000000_000000000_010001010_001000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000011_011111110_001100011_000000000_000000000_000000000_000000000_010111101_010001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011111110_001101011_000000000_000000000_000000000_001010101_011100101_001011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_011000100_011100100_000001011_000000000_000000000_010011010_011111110_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011111110_010000001_000000001_000001001_011001111_011111111_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000001_011111110_010110111_010111100_010101111_011111110_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_001110100_010010011_000010110_010010010_011111110_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111110_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111110_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100111_011111110_000111001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010000111_011101000_000001000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011111011_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100011_011110110_000101001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111110_011100101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_97 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101101_010011010_011010000_011111000_011100110_011111110_011111111_010001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_011001101_011111110_011111110_011111110_011111110_011111110_011111110_011010101_000011111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011010010_011111110_011111110_011111110_011111110_011101100_011111110_011111110_011111110_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100010_011111110_011111110_011111110_010011000_000101000_000011010_010010111_011111110_011111110_010101000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100110_011111110_011111110_011001010_000101100_000000000_000001010_011001111_011111110_011111110_011001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110101_011111100_011111110_011110010_001010011_010001000_010110100_011111110_011111110_011111110_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010111101_011111110_011111110_011111110_011111110_011111110_011111110_011111110_011111110_000111111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_000111000_011010001_011111110_011111110_011111110_011111110_011111110_011001001_000000001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011100100_011111110_011111110_011111110_011101110_001011100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100111_011111000_011111110_011111110_011111110_000111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_011111000_011111110_011111110_011111101_010100110_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001100100_011100110_011111110_011111110_010101010_001110001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011111101_011111110_011111110_011100101_000010000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011111_011100011_011111110_011111110_011111110_010000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100110_011100100_011111110_011111110_011111110_011001010_000010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011000001_011111110_011111110_011111110_011001010_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011011_011110110_011111110_011111110_011110010_001011010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000100011_011110010_011111110_011111110_011111110_010001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010110_011111110_011111110_010111001_000010111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010110111_011111110_011110111_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_98 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000110_011001010_011111111_001111110_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011101111_011111101_011111101_011111101_000001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010001_011110010_011111101_011000001_010100110_011111101_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110100_011001010_011111101_010110100_000000111_000111100_011111101_001110111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001001000_011010011_011111000_001100111_000001110_000000000_000111100_011111101_010011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000010_011110100_011111010_010000110_000000000_000001001_001111011_011101001_011111101_010101111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000010000_011101000_011111101_010010010_000110100_010011101_011101001_011111101_011111101_011111101_000110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110110_011110101_011111101_011010000_011111001_011111101_011111101_011111101_011111101_011011100_000000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011011100_011111101_011111101_011110000_011111101_011111101_011111100_010111010_000001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_001011100_001011100_000101111_011111101_011111101_010001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010100100_011111101_010001101_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010010_011111100_011111101_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011110_011111101_011011001_000010010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101000_011110010_011110111_001001101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010011001_011111101_011100010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001000_011011111_011111101_001100110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001011_011111101_011111101_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110110_011111101_011111101_000111010_001110110_000110110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101011_011111101_011111101_011111101_011101110_000100111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_010101011_011111101_011001000_001000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
parameter data_99 = 7056'b000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000110_001110100_011110011_011100000_011110110_000111011_000000000_000011111_001111001_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000010_010010101_010111111_001011111_000001000_010011110_000011001_000010001_011011011_011100100_000010101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000001110_010101101_010010101_000111000_000000000_000000000_000111101_000000101_011000110_011100100_000101100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001010110_011001000_000011001_000000000_000000000_000000000_000000000_001000010_011001011_001001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001111101_010001010_000000000_000000000_000000000_000000000_000101011_011110011_011100110_000101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_010001011_011001001_000000110_000000000_000000000_000000000_000000000_010010101_011111100_001010100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011000_011100100_000001010_000000000_000000000_000000000_000010010_010011000_011111101_010001011_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000100_011100001_001100000_000000000_000000000_000000010_001000100_011000010_011100000_001101110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000110001_011100101_000010100_000011100_000111100_010010111_011111111_011111001_001000111_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000101001_011111001_011001110_011111101_011011101_011001110_011110110_011001010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101010_011000100_001111011_000010000_010000111_011110110_010001110_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001101110_011111110_011000110_000000101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011101_011111010_011101101_000011001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000011_011011011_011010010_000011000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001110000_011110100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001000000_011110100_001111100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_001011110_011101001_010100100_000000100_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_011011110_000001001_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_011010011_001111101_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000011000_001011010_000000010_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000_000000000;
